
module up_counter_WIDTH14_1_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
endmodule


module up_counter_WIDTH14_1 ( clk, rst, clr, count, en_BAR );
  output [13:0] count;
  input clk, rst, clr, en_BAR;
  wire   en, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n1, n2,
         n3, n4;
  assign en = en_BAR;

  up_counter_WIDTH14_1_DW01_inc_0 add_18 ( .A(count), .SUM({N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  DFFRX1 \count_reg[5]  ( .D(n13), .CK(clk), .RN(n3), .Q(count[5]) );
  DFFRX1 \count_reg[4]  ( .D(n14), .CK(clk), .RN(n3), .Q(count[4]) );
  DFFRX1 \count_reg[3]  ( .D(n15), .CK(clk), .RN(n3), .Q(count[3]) );
  DFFRX1 \count_reg[2]  ( .D(n16), .CK(clk), .RN(n3), .Q(count[2]) );
  DFFRX1 \count_reg[1]  ( .D(n17), .CK(clk), .RN(n3), .Q(count[1]) );
  DFFRX1 \count_reg[0]  ( .D(n2), .CK(clk), .RN(n3), .Q(count[0]) );
  DFFRX1 \count_reg[6]  ( .D(n12), .CK(clk), .RN(n3), .Q(count[6]) );
  DFFRX1 \count_reg[7]  ( .D(n11), .CK(clk), .RN(n3), .Q(count[7]) );
  DFFRX1 \count_reg[8]  ( .D(n10), .CK(clk), .RN(n3), .Q(count[8]) );
  DFFRX1 \count_reg[9]  ( .D(n9), .CK(clk), .RN(n3), .Q(count[9]) );
  DFFRX1 \count_reg[10]  ( .D(n8), .CK(clk), .RN(n3), .Q(count[10]) );
  DFFRX1 \count_reg[11]  ( .D(n7), .CK(clk), .RN(n3), .Q(count[11]) );
  DFFRX1 \count_reg[12]  ( .D(n6), .CK(clk), .RN(n3), .Q(count[12]) );
  DFFRX1 \count_reg[13]  ( .D(n5), .CK(clk), .RN(n3), .Q(count[13]) );
  INVX3 U3 ( .A(en), .Y(n1) );
  AO22X1 U4 ( .A0(N4), .A1(n1), .B0(count[0]), .B1(n4), .Y(n2) );
  INVX3 U5 ( .A(n1), .Y(n4) );
  INVX3 U6 ( .A(rst), .Y(n3) );
  AO22X1 U7 ( .A0(count[13]), .A1(n4), .B0(N17), .B1(n1), .Y(n5) );
  AO22X1 U8 ( .A0(count[12]), .A1(n4), .B0(N16), .B1(n1), .Y(n6) );
  AO22X1 U9 ( .A0(count[11]), .A1(n4), .B0(N15), .B1(n1), .Y(n7) );
  AO22X1 U10 ( .A0(count[10]), .A1(n4), .B0(N14), .B1(n1), .Y(n8) );
  AO22X1 U11 ( .A0(count[9]), .A1(n4), .B0(N13), .B1(n1), .Y(n9) );
  AO22X1 U12 ( .A0(count[8]), .A1(n4), .B0(N12), .B1(n1), .Y(n10) );
  AO22X1 U13 ( .A0(count[7]), .A1(n4), .B0(N11), .B1(n1), .Y(n11) );
  AO22X1 U14 ( .A0(count[6]), .A1(n4), .B0(N10), .B1(n1), .Y(n12) );
  AO22X1 U15 ( .A0(count[5]), .A1(n4), .B0(N9), .B1(n1), .Y(n13) );
  AO22X1 U16 ( .A0(count[4]), .A1(n4), .B0(N8), .B1(n1), .Y(n14) );
  AO22X1 U17 ( .A0(count[3]), .A1(n4), .B0(N7), .B1(n1), .Y(n15) );
  AO22X1 U18 ( .A0(count[2]), .A1(n4), .B0(N6), .B1(n1), .Y(n16) );
  AO22X1 U19 ( .A0(count[1]), .A1(n4), .B0(N5), .B1(n1), .Y(n17) );
endmodule


module up_counter_WIDTH14_0_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
endmodule


module up_counter_WIDTH14_0 ( clk, rst, en, clr, count );
  output [13:0] count;
  input clk, rst, en, clr;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, n1,
         n2, n3, n4, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30;

  up_counter_WIDTH14_0_DW01_inc_0 add_18 ( .A(count), .SUM({N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  DFFRX1 \count_reg[2]  ( .D(n19), .CK(clk), .RN(n3), .Q(count[2]) );
  DFFRX1 \count_reg[1]  ( .D(n18), .CK(clk), .RN(n3), .Q(count[1]) );
  DFFRX1 \count_reg[0]  ( .D(n1), .CK(clk), .RN(n3), .Q(count[0]) );
  DFFRX1 \count_reg[3]  ( .D(n20), .CK(clk), .RN(n3), .Q(count[3]) );
  DFFRX1 \count_reg[4]  ( .D(n21), .CK(clk), .RN(n3), .Q(count[4]) );
  DFFRX1 \count_reg[5]  ( .D(n22), .CK(clk), .RN(n3), .Q(count[5]) );
  DFFRX1 \count_reg[6]  ( .D(n23), .CK(clk), .RN(n3), .Q(count[6]) );
  DFFRX1 \count_reg[7]  ( .D(n24), .CK(clk), .RN(n3), .Q(count[7]) );
  DFFRX1 \count_reg[8]  ( .D(n25), .CK(clk), .RN(n3), .Q(count[8]) );
  DFFRX1 \count_reg[9]  ( .D(n26), .CK(clk), .RN(n3), .Q(count[9]) );
  DFFRX1 \count_reg[10]  ( .D(n27), .CK(clk), .RN(n3), .Q(count[10]) );
  DFFRX1 \count_reg[11]  ( .D(n28), .CK(clk), .RN(n3), .Q(count[11]) );
  DFFRX1 \count_reg[12]  ( .D(n29), .CK(clk), .RN(n3), .Q(count[12]) );
  DFFRX1 \count_reg[13]  ( .D(n30), .CK(clk), .RN(n3), .Q(count[13]) );
  AO22X1 U3 ( .A0(N4), .A1(n2), .B0(count[0]), .B1(n4), .Y(n1) );
  INVX3 U4 ( .A(n2), .Y(n4) );
  INVX3 U5 ( .A(rst), .Y(n3) );
  AO22X1 U6 ( .A0(count[13]), .A1(n4), .B0(N17), .B1(n2), .Y(n30) );
  AO22X1 U7 ( .A0(count[12]), .A1(n4), .B0(N16), .B1(n2), .Y(n29) );
  AO22X1 U8 ( .A0(count[11]), .A1(n4), .B0(N15), .B1(n2), .Y(n28) );
  AO22X1 U9 ( .A0(count[10]), .A1(n4), .B0(N14), .B1(n2), .Y(n27) );
  AO22X1 U10 ( .A0(count[9]), .A1(n4), .B0(N13), .B1(n2), .Y(n26) );
  AO22X1 U11 ( .A0(count[8]), .A1(n4), .B0(N12), .B1(n2), .Y(n25) );
  AO22X1 U12 ( .A0(count[7]), .A1(n4), .B0(N11), .B1(n2), .Y(n24) );
  CLKBUFX3 U13 ( .A(en), .Y(n2) );
  AO22X1 U14 ( .A0(count[6]), .A1(n4), .B0(N10), .B1(n2), .Y(n23) );
  AO22X1 U15 ( .A0(count[5]), .A1(n4), .B0(N9), .B1(n2), .Y(n22) );
  AO22X1 U16 ( .A0(count[4]), .A1(n4), .B0(N8), .B1(n2), .Y(n21) );
  AO22X1 U17 ( .A0(count[3]), .A1(n4), .B0(N7), .B1(n2), .Y(n20) );
  AO22X1 U18 ( .A0(count[2]), .A1(n4), .B0(N6), .B1(n2), .Y(n19) );
  AO22X1 U19 ( .A0(count[1]), .A1(n4), .B0(N5), .B1(n2), .Y(n18) );
endmodule


module up_counter_WIDTH7_1_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module up_counter_WIDTH7_1 ( clk, rst, en, clr, count );
  output [6:0] count;
  input clk, rst, en, clr;
  wire   N4, N5, N6, N7, N8, N9, N10, n5, n6, n7, n8, n9, n10, n1, n2, n3;

  up_counter_WIDTH7_1_DW01_inc_0 add_18 ( .A(count), .SUM({N10, N9, N8, N7, N6, 
        N5, N4}) );
  DFFRX2 \count_reg[0]  ( .D(n1), .CK(clk), .RN(n3), .Q(count[0]) );
  DFFRX2 \count_reg[5]  ( .D(n6), .CK(clk), .RN(n3), .Q(count[5]) );
  DFFRX2 \count_reg[4]  ( .D(n7), .CK(clk), .RN(n3), .Q(count[4]) );
  DFFRX1 \count_reg[3]  ( .D(n8), .CK(clk), .RN(n3), .Q(count[3]) );
  DFFRX1 \count_reg[2]  ( .D(n9), .CK(clk), .RN(n3), .Q(count[2]) );
  DFFRX1 \count_reg[1]  ( .D(n10), .CK(clk), .RN(n3), .Q(count[1]) );
  DFFRHQX2 \count_reg[6]  ( .D(n5), .CK(clk), .RN(n3), .Q(count[6]) );
  AO22X1 U3 ( .A0(N4), .A1(en), .B0(count[0]), .B1(n2), .Y(n1) );
  CLKINVX1 U4 ( .A(en), .Y(n2) );
  INVX3 U5 ( .A(rst), .Y(n3) );
  AO22X1 U6 ( .A0(count[6]), .A1(n2), .B0(N10), .B1(en), .Y(n5) );
  AO22XL U7 ( .A0(count[4]), .A1(n2), .B0(N8), .B1(en), .Y(n7) );
  AO22X1 U8 ( .A0(count[5]), .A1(n2), .B0(N9), .B1(en), .Y(n6) );
  AO22X1 U9 ( .A0(count[3]), .A1(n2), .B0(N7), .B1(en), .Y(n8) );
  AO22X1 U10 ( .A0(count[1]), .A1(n2), .B0(N5), .B1(en), .Y(n10) );
  AO22X1 U11 ( .A0(count[2]), .A1(n2), .B0(N6), .B1(en), .Y(n9) );
endmodule


module line_buffer_1_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVXL U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module line_buffer_1 ( clk, rst, en, data_in, data_out, valid );
  input [7:0] data_in;
  output [7:0] data_out;
  input clk, rst, en;
  output valid;
  wire   N26, N27, N28, N29, N30, N31, N32, \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] ,
         \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] ,
         \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] ,
         \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] ,
         \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] ,
         \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[15][7] , \mem[15][6] ,
         \mem[15][5] , \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] ,
         \mem[15][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] , \mem[16][4] ,
         \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] ,
         \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] ,
         \mem[19][7] , \mem[19][6] , \mem[19][5] , \mem[19][4] , \mem[19][3] ,
         \mem[19][2] , \mem[19][1] , \mem[19][0] , \mem[20][7] , \mem[20][6] ,
         \mem[20][5] , \mem[20][4] , \mem[20][3] , \mem[20][2] , \mem[20][1] ,
         \mem[20][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] , \mem[21][4] ,
         \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] ,
         \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] ,
         \mem[24][7] , \mem[24][6] , \mem[24][5] , \mem[24][4] , \mem[24][3] ,
         \mem[24][2] , \mem[24][1] , \mem[24][0] , \mem[25][7] , \mem[25][6] ,
         \mem[25][5] , \mem[25][4] , \mem[25][3] , \mem[25][2] , \mem[25][1] ,
         \mem[25][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] , \mem[26][4] ,
         \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] ,
         \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] ,
         \mem[29][7] , \mem[29][6] , \mem[29][5] , \mem[29][4] , \mem[29][3] ,
         \mem[29][2] , \mem[29][1] , \mem[29][0] , \mem[30][7] , \mem[30][6] ,
         \mem[30][5] , \mem[30][4] , \mem[30][3] , \mem[30][2] , \mem[30][1] ,
         \mem[30][0] , \mem[31][7] , \mem[31][6] , \mem[31][5] , \mem[31][4] ,
         \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] , \mem[32][7] ,
         \mem[32][6] , \mem[32][5] , \mem[32][4] , \mem[32][3] , \mem[32][2] ,
         \mem[32][1] , \mem[32][0] , \mem[33][7] , \mem[33][6] , \mem[33][5] ,
         \mem[33][4] , \mem[33][3] , \mem[33][2] , \mem[33][1] , \mem[33][0] ,
         \mem[34][7] , \mem[34][6] , \mem[34][5] , \mem[34][4] , \mem[34][3] ,
         \mem[34][2] , \mem[34][1] , \mem[34][0] , \mem[35][7] , \mem[35][6] ,
         \mem[35][5] , \mem[35][4] , \mem[35][3] , \mem[35][2] , \mem[35][1] ,
         \mem[35][0] , \mem[36][7] , \mem[36][6] , \mem[36][5] , \mem[36][4] ,
         \mem[36][3] , \mem[36][2] , \mem[36][1] , \mem[36][0] , \mem[37][7] ,
         \mem[37][6] , \mem[37][5] , \mem[37][4] , \mem[37][3] , \mem[37][2] ,
         \mem[37][1] , \mem[37][0] , \mem[38][7] , \mem[38][6] , \mem[38][5] ,
         \mem[38][4] , \mem[38][3] , \mem[38][2] , \mem[38][1] , \mem[38][0] ,
         \mem[39][7] , \mem[39][6] , \mem[39][5] , \mem[39][4] , \mem[39][3] ,
         \mem[39][2] , \mem[39][1] , \mem[39][0] , \mem[40][7] , \mem[40][6] ,
         \mem[40][5] , \mem[40][4] , \mem[40][3] , \mem[40][2] , \mem[40][1] ,
         \mem[40][0] , \mem[41][7] , \mem[41][6] , \mem[41][5] , \mem[41][4] ,
         \mem[41][3] , \mem[41][2] , \mem[41][1] , \mem[41][0] , \mem[42][7] ,
         \mem[42][6] , \mem[42][5] , \mem[42][4] , \mem[42][3] , \mem[42][2] ,
         \mem[42][1] , \mem[42][0] , \mem[43][7] , \mem[43][6] , \mem[43][5] ,
         \mem[43][4] , \mem[43][3] , \mem[43][2] , \mem[43][1] , \mem[43][0] ,
         \mem[44][7] , \mem[44][6] , \mem[44][5] , \mem[44][4] , \mem[44][3] ,
         \mem[44][2] , \mem[44][1] , \mem[44][0] , \mem[45][7] , \mem[45][6] ,
         \mem[45][5] , \mem[45][4] , \mem[45][3] , \mem[45][2] , \mem[45][1] ,
         \mem[45][0] , \mem[46][7] , \mem[46][6] , \mem[46][5] , \mem[46][4] ,
         \mem[46][3] , \mem[46][2] , \mem[46][1] , \mem[46][0] , \mem[47][7] ,
         \mem[47][6] , \mem[47][5] , \mem[47][4] , \mem[47][3] , \mem[47][2] ,
         \mem[47][1] , \mem[47][0] , \mem[48][7] , \mem[48][6] , \mem[48][5] ,
         \mem[48][4] , \mem[48][3] , \mem[48][2] , \mem[48][1] , \mem[48][0] ,
         \mem[49][7] , \mem[49][6] , \mem[49][5] , \mem[49][4] , \mem[49][3] ,
         \mem[49][2] , \mem[49][1] , \mem[49][0] , \mem[50][7] , \mem[50][6] ,
         \mem[50][5] , \mem[50][4] , \mem[50][3] , \mem[50][2] , \mem[50][1] ,
         \mem[50][0] , \mem[51][7] , \mem[51][6] , \mem[51][5] , \mem[51][4] ,
         \mem[51][3] , \mem[51][2] , \mem[51][1] , \mem[51][0] , \mem[52][7] ,
         \mem[52][6] , \mem[52][5] , \mem[52][4] , \mem[52][3] , \mem[52][2] ,
         \mem[52][1] , \mem[52][0] , \mem[53][7] , \mem[53][6] , \mem[53][5] ,
         \mem[53][4] , \mem[53][3] , \mem[53][2] , \mem[53][1] , \mem[53][0] ,
         \mem[54][7] , \mem[54][6] , \mem[54][5] , \mem[54][4] , \mem[54][3] ,
         \mem[54][2] , \mem[54][1] , \mem[54][0] , \mem[55][7] , \mem[55][6] ,
         \mem[55][5] , \mem[55][4] , \mem[55][3] , \mem[55][2] , \mem[55][1] ,
         \mem[55][0] , \mem[56][7] , \mem[56][6] , \mem[56][5] , \mem[56][4] ,
         \mem[56][3] , \mem[56][2] , \mem[56][1] , \mem[56][0] , \mem[57][7] ,
         \mem[57][6] , \mem[57][5] , \mem[57][4] , \mem[57][3] , \mem[57][2] ,
         \mem[57][1] , \mem[57][0] , \mem[58][7] , \mem[58][6] , \mem[58][5] ,
         \mem[58][4] , \mem[58][3] , \mem[58][2] , \mem[58][1] , \mem[58][0] ,
         \mem[59][7] , \mem[59][6] , \mem[59][5] , \mem[59][4] , \mem[59][3] ,
         \mem[59][2] , \mem[59][1] , \mem[59][0] , \mem[60][7] , \mem[60][6] ,
         \mem[60][5] , \mem[60][4] , \mem[60][3] , \mem[60][2] , \mem[60][1] ,
         \mem[60][0] , \mem[61][7] , \mem[61][6] , \mem[61][5] , \mem[61][4] ,
         \mem[61][3] , \mem[61][2] , \mem[61][1] , \mem[61][0] , \mem[62][7] ,
         \mem[62][6] , \mem[62][5] , \mem[62][4] , \mem[62][3] , \mem[62][2] ,
         \mem[62][1] , \mem[62][0] , \mem[63][7] , \mem[63][6] , \mem[63][5] ,
         \mem[63][4] , \mem[63][3] , \mem[63][2] , \mem[63][1] , \mem[63][0] ,
         \mem[64][7] , \mem[64][6] , \mem[64][5] , \mem[64][4] , \mem[64][3] ,
         \mem[64][2] , \mem[64][1] , \mem[64][0] , \mem[65][7] , \mem[65][6] ,
         \mem[65][5] , \mem[65][4] , \mem[65][3] , \mem[65][2] , \mem[65][1] ,
         \mem[65][0] , \mem[66][7] , \mem[66][6] , \mem[66][5] , \mem[66][4] ,
         \mem[66][3] , \mem[66][2] , \mem[66][1] , \mem[66][0] , \mem[67][7] ,
         \mem[67][6] , \mem[67][5] , \mem[67][4] , \mem[67][3] , \mem[67][2] ,
         \mem[67][1] , \mem[67][0] , \mem[68][7] , \mem[68][6] , \mem[68][5] ,
         \mem[68][4] , \mem[68][3] , \mem[68][2] , \mem[68][1] , \mem[68][0] ,
         \mem[69][7] , \mem[69][6] , \mem[69][5] , \mem[69][4] , \mem[69][3] ,
         \mem[69][2] , \mem[69][1] , \mem[69][0] , \mem[70][7] , \mem[70][6] ,
         \mem[70][5] , \mem[70][4] , \mem[70][3] , \mem[70][2] , \mem[70][1] ,
         \mem[70][0] , \mem[71][7] , \mem[71][6] , \mem[71][5] , \mem[71][4] ,
         \mem[71][3] , \mem[71][2] , \mem[71][1] , \mem[71][0] , \mem[72][7] ,
         \mem[72][6] , \mem[72][5] , \mem[72][4] , \mem[72][3] , \mem[72][2] ,
         \mem[72][1] , \mem[72][0] , \mem[73][7] , \mem[73][6] , \mem[73][5] ,
         \mem[73][4] , \mem[73][3] , \mem[73][2] , \mem[73][1] , \mem[73][0] ,
         \mem[74][7] , \mem[74][6] , \mem[74][5] , \mem[74][4] , \mem[74][3] ,
         \mem[74][2] , \mem[74][1] , \mem[74][0] , \mem[75][7] , \mem[75][6] ,
         \mem[75][5] , \mem[75][4] , \mem[75][3] , \mem[75][2] , \mem[75][1] ,
         \mem[75][0] , \mem[76][7] , \mem[76][6] , \mem[76][5] , \mem[76][4] ,
         \mem[76][3] , \mem[76][2] , \mem[76][1] , \mem[76][0] , \mem[77][7] ,
         \mem[77][6] , \mem[77][5] , \mem[77][4] , \mem[77][3] , \mem[77][2] ,
         \mem[77][1] , \mem[77][0] , \mem[78][7] , \mem[78][6] , \mem[78][5] ,
         \mem[78][4] , \mem[78][3] , \mem[78][2] , \mem[78][1] , \mem[78][0] ,
         \mem[79][7] , \mem[79][6] , \mem[79][5] , \mem[79][4] , \mem[79][3] ,
         \mem[79][2] , \mem[79][1] , \mem[79][0] , \mem[80][7] , \mem[80][6] ,
         \mem[80][5] , \mem[80][4] , \mem[80][3] , \mem[80][2] , \mem[80][1] ,
         \mem[80][0] , \mem[81][7] , \mem[81][6] , \mem[81][5] , \mem[81][4] ,
         \mem[81][3] , \mem[81][2] , \mem[81][1] , \mem[81][0] , \mem[82][7] ,
         \mem[82][6] , \mem[82][5] , \mem[82][4] , \mem[82][3] , \mem[82][2] ,
         \mem[82][1] , \mem[82][0] , \mem[83][7] , \mem[83][6] , \mem[83][5] ,
         \mem[83][4] , \mem[83][3] , \mem[83][2] , \mem[83][1] , \mem[83][0] ,
         \mem[84][7] , \mem[84][6] , \mem[84][5] , \mem[84][4] , \mem[84][3] ,
         \mem[84][2] , \mem[84][1] , \mem[84][0] , \mem[85][7] , \mem[85][6] ,
         \mem[85][5] , \mem[85][4] , \mem[85][3] , \mem[85][2] , \mem[85][1] ,
         \mem[85][0] , \mem[86][7] , \mem[86][6] , \mem[86][5] , \mem[86][4] ,
         \mem[86][3] , \mem[86][2] , \mem[86][1] , \mem[86][0] , \mem[87][7] ,
         \mem[87][6] , \mem[87][5] , \mem[87][4] , \mem[87][3] , \mem[87][2] ,
         \mem[87][1] , \mem[87][0] , \mem[88][7] , \mem[88][6] , \mem[88][5] ,
         \mem[88][4] , \mem[88][3] , \mem[88][2] , \mem[88][1] , \mem[88][0] ,
         \mem[89][7] , \mem[89][6] , \mem[89][5] , \mem[89][4] , \mem[89][3] ,
         \mem[89][2] , \mem[89][1] , \mem[89][0] , \mem[90][7] , \mem[90][6] ,
         \mem[90][5] , \mem[90][4] , \mem[90][3] , \mem[90][2] , \mem[90][1] ,
         \mem[90][0] , \mem[91][7] , \mem[91][6] , \mem[91][5] , \mem[91][4] ,
         \mem[91][3] , \mem[91][2] , \mem[91][1] , \mem[91][0] , \mem[92][7] ,
         \mem[92][6] , \mem[92][5] , \mem[92][4] , \mem[92][3] , \mem[92][2] ,
         \mem[92][1] , \mem[92][0] , \mem[93][7] , \mem[93][6] , \mem[93][5] ,
         \mem[93][4] , \mem[93][3] , \mem[93][2] , \mem[93][1] , \mem[93][0] ,
         \mem[94][7] , \mem[94][6] , \mem[94][5] , \mem[94][4] , \mem[94][3] ,
         \mem[94][2] , \mem[94][1] , \mem[94][0] , \mem[95][7] , \mem[95][6] ,
         \mem[95][5] , \mem[95][4] , \mem[95][3] , \mem[95][2] , \mem[95][1] ,
         \mem[95][0] , \mem[96][7] , \mem[96][6] , \mem[96][5] , \mem[96][4] ,
         \mem[96][3] , \mem[96][2] , \mem[96][1] , \mem[96][0] , \mem[97][7] ,
         \mem[97][6] , \mem[97][5] , \mem[97][4] , \mem[97][3] , \mem[97][2] ,
         \mem[97][1] , \mem[97][0] , \mem[98][7] , \mem[98][6] , \mem[98][5] ,
         \mem[98][4] , \mem[98][3] , \mem[98][2] , \mem[98][1] , \mem[98][0] ,
         \mem[99][7] , \mem[99][6] , \mem[99][5] , \mem[99][4] , \mem[99][3] ,
         \mem[99][2] , \mem[99][1] , \mem[99][0] , \mem[100][7] ,
         \mem[100][6] , \mem[100][5] , \mem[100][4] , \mem[100][3] ,
         \mem[100][2] , \mem[100][1] , \mem[100][0] , \mem[101][7] ,
         \mem[101][6] , \mem[101][5] , \mem[101][4] , \mem[101][3] ,
         \mem[101][2] , \mem[101][1] , \mem[101][0] , \mem[102][7] ,
         \mem[102][6] , \mem[102][5] , \mem[102][4] , \mem[102][3] ,
         \mem[102][2] , \mem[102][1] , \mem[102][0] , \mem[103][7] ,
         \mem[103][6] , \mem[103][5] , \mem[103][4] , \mem[103][3] ,
         \mem[103][2] , \mem[103][1] , \mem[103][0] , \mem[104][7] ,
         \mem[104][6] , \mem[104][5] , \mem[104][4] , \mem[104][3] ,
         \mem[104][2] , \mem[104][1] , \mem[104][0] , \mem[105][7] ,
         \mem[105][6] , \mem[105][5] , \mem[105][4] , \mem[105][3] ,
         \mem[105][2] , \mem[105][1] , \mem[105][0] , \mem[106][7] ,
         \mem[106][6] , \mem[106][5] , \mem[106][4] , \mem[106][3] ,
         \mem[106][2] , \mem[106][1] , \mem[106][0] , \mem[107][7] ,
         \mem[107][6] , \mem[107][5] , \mem[107][4] , \mem[107][3] ,
         \mem[107][2] , \mem[107][1] , \mem[107][0] , \mem[108][7] ,
         \mem[108][6] , \mem[108][5] , \mem[108][4] , \mem[108][3] ,
         \mem[108][2] , \mem[108][1] , \mem[108][0] , \mem[109][7] ,
         \mem[109][6] , \mem[109][5] , \mem[109][4] , \mem[109][3] ,
         \mem[109][2] , \mem[109][1] , \mem[109][0] , \mem[110][7] ,
         \mem[110][6] , \mem[110][5] , \mem[110][4] , \mem[110][3] ,
         \mem[110][2] , \mem[110][1] , \mem[110][0] , \mem[111][7] ,
         \mem[111][6] , \mem[111][5] , \mem[111][4] , \mem[111][3] ,
         \mem[111][2] , \mem[111][1] , \mem[111][0] , \mem[112][7] ,
         \mem[112][6] , \mem[112][5] , \mem[112][4] , \mem[112][3] ,
         \mem[112][2] , \mem[112][1] , \mem[112][0] , \mem[113][7] ,
         \mem[113][6] , \mem[113][5] , \mem[113][4] , \mem[113][3] ,
         \mem[113][2] , \mem[113][1] , \mem[113][0] , \mem[114][7] ,
         \mem[114][6] , \mem[114][5] , \mem[114][4] , \mem[114][3] ,
         \mem[114][2] , \mem[114][1] , \mem[114][0] , \mem[115][7] ,
         \mem[115][6] , \mem[115][5] , \mem[115][4] , \mem[115][3] ,
         \mem[115][2] , \mem[115][1] , \mem[115][0] , \mem[116][7] ,
         \mem[116][6] , \mem[116][5] , \mem[116][4] , \mem[116][3] ,
         \mem[116][2] , \mem[116][1] , \mem[116][0] , \mem[117][7] ,
         \mem[117][6] , \mem[117][5] , \mem[117][4] , \mem[117][3] ,
         \mem[117][2] , \mem[117][1] , \mem[117][0] , \mem[118][7] ,
         \mem[118][6] , \mem[118][5] , \mem[118][4] , \mem[118][3] ,
         \mem[118][2] , \mem[118][1] , \mem[118][0] , \mem[119][7] ,
         \mem[119][6] , \mem[119][5] , \mem[119][4] , \mem[119][3] ,
         \mem[119][2] , \mem[119][1] , \mem[119][0] , \mem[120][7] ,
         \mem[120][6] , \mem[120][5] , \mem[120][4] , \mem[120][3] ,
         \mem[120][2] , \mem[120][1] , \mem[120][0] , \mem[121][7] ,
         \mem[121][6] , \mem[121][5] , \mem[121][4] , \mem[121][3] ,
         \mem[121][2] , \mem[121][1] , \mem[121][0] , \mem[122][7] ,
         \mem[122][6] , \mem[122][5] , \mem[122][4] , \mem[122][3] ,
         \mem[122][2] , \mem[122][1] , \mem[122][0] , \mem[123][7] ,
         \mem[123][6] , \mem[123][5] , \mem[123][4] , \mem[123][3] ,
         \mem[123][2] , \mem[123][1] , \mem[123][0] , \mem[124][7] ,
         \mem[124][6] , \mem[124][5] , \mem[124][4] , \mem[124][3] ,
         \mem[124][2] , \mem[124][1] , \mem[124][0] , \mem[125][7] ,
         \mem[125][6] , \mem[125][5] , \mem[125][4] , \mem[125][3] ,
         \mem[125][2] , \mem[125][1] , \mem[125][0] , \mem[126][7] ,
         \mem[126][6] , \mem[126][5] , \mem[126][4] , \mem[126][3] ,
         \mem[126][2] , \mem[126][1] , \mem[126][0] , \mem[127][7] ,
         \mem[127][6] , \mem[127][5] , \mem[127][4] , \mem[127][3] ,
         \mem[127][2] , \mem[127][1] , \mem[127][0] , N33, N34, N35, N36, N37,
         N38, N39, N40, N41, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n435,
         n436, n437, n438, n439, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062;
  wire   [6:0] write_counter_count;
  wire   [0:127] valid_mem;

  up_counter_WIDTH7_1 write_counter ( .clk(clk), .rst(rst), .en(n912), .clr(
        1'b0), .count(write_counter_count) );
  line_buffer_1_DW01_inc_0 add_15 ( .A(write_counter_count), .SUM({N32, N31, 
        N30, N29, N28, N27, N26}) );
  EDFFX1 \mem_reg[1][7]  ( .D(n911), .E(n956), .CK(clk), .Q(\mem[1][7] ) );
  EDFFX1 \mem_reg[1][6]  ( .D(n906), .E(n956), .CK(clk), .Q(\mem[1][6] ) );
  EDFFX1 \mem_reg[1][5]  ( .D(n901), .E(n956), .CK(clk), .Q(\mem[1][5] ) );
  EDFFX1 \mem_reg[1][4]  ( .D(n896), .E(n956), .CK(clk), .Q(\mem[1][4] ) );
  EDFFX1 \mem_reg[1][3]  ( .D(n891), .E(n956), .CK(clk), .Q(\mem[1][3] ) );
  EDFFX1 \mem_reg[1][2]  ( .D(n886), .E(n956), .CK(clk), .Q(\mem[1][2] ) );
  EDFFX1 \mem_reg[1][1]  ( .D(n881), .E(n956), .CK(clk), .Q(\mem[1][1] ) );
  EDFFX1 \mem_reg[1][0]  ( .D(n876), .E(n956), .CK(clk), .Q(\mem[1][0] ) );
  EDFFX1 \mem_reg[5][7]  ( .D(n911), .E(n965), .CK(clk), .Q(\mem[5][7] ) );
  EDFFX1 \mem_reg[5][6]  ( .D(n906), .E(n965), .CK(clk), .Q(\mem[5][6] ) );
  EDFFX1 \mem_reg[5][5]  ( .D(n901), .E(n965), .CK(clk), .Q(\mem[5][5] ) );
  EDFFX1 \mem_reg[5][4]  ( .D(n896), .E(n965), .CK(clk), .Q(\mem[5][4] ) );
  EDFFX1 \mem_reg[5][3]  ( .D(n891), .E(n965), .CK(clk), .Q(\mem[5][3] ) );
  EDFFX1 \mem_reg[5][2]  ( .D(n886), .E(n965), .CK(clk), .Q(\mem[5][2] ) );
  EDFFX1 \mem_reg[5][1]  ( .D(n881), .E(n965), .CK(clk), .Q(\mem[5][1] ) );
  EDFFX1 \mem_reg[5][0]  ( .D(n876), .E(n965), .CK(clk), .Q(\mem[5][0] ) );
  EDFFX1 \mem_reg[9][7]  ( .D(n908), .E(n974), .CK(clk), .Q(\mem[9][7] ) );
  EDFFX1 \mem_reg[9][6]  ( .D(n903), .E(n974), .CK(clk), .Q(\mem[9][6] ) );
  EDFFX1 \mem_reg[9][5]  ( .D(n898), .E(n974), .CK(clk), .Q(\mem[9][5] ) );
  EDFFX1 \mem_reg[9][4]  ( .D(n893), .E(n974), .CK(clk), .Q(\mem[9][4] ) );
  EDFFX1 \mem_reg[9][3]  ( .D(n888), .E(n974), .CK(clk), .Q(\mem[9][3] ) );
  EDFFX1 \mem_reg[9][2]  ( .D(n883), .E(n974), .CK(clk), .Q(\mem[9][2] ) );
  EDFFX1 \mem_reg[9][1]  ( .D(n878), .E(n974), .CK(clk), .Q(\mem[9][1] ) );
  EDFFX1 \mem_reg[9][0]  ( .D(n873), .E(n974), .CK(clk), .Q(\mem[9][0] ) );
  EDFFX1 \mem_reg[13][7]  ( .D(n907), .E(n983), .CK(clk), .Q(\mem[13][7] ) );
  EDFFX1 \mem_reg[13][6]  ( .D(n902), .E(n983), .CK(clk), .Q(\mem[13][6] ) );
  EDFFX1 \mem_reg[13][5]  ( .D(n897), .E(n983), .CK(clk), .Q(\mem[13][5] ) );
  EDFFX1 \mem_reg[13][4]  ( .D(n892), .E(n983), .CK(clk), .Q(\mem[13][4] ) );
  EDFFX1 \mem_reg[13][3]  ( .D(n887), .E(n983), .CK(clk), .Q(\mem[13][3] ) );
  EDFFX1 \mem_reg[13][2]  ( .D(n882), .E(n983), .CK(clk), .Q(\mem[13][2] ) );
  EDFFX1 \mem_reg[13][1]  ( .D(n877), .E(n983), .CK(clk), .Q(\mem[13][1] ) );
  EDFFX1 \mem_reg[13][0]  ( .D(n872), .E(n983), .CK(clk), .Q(\mem[13][0] ) );
  EDFFX1 \mem_reg[17][7]  ( .D(n909), .E(n955), .CK(clk), .Q(\mem[17][7] ) );
  EDFFX1 \mem_reg[17][6]  ( .D(n904), .E(n955), .CK(clk), .Q(\mem[17][6] ) );
  EDFFX1 \mem_reg[17][5]  ( .D(n899), .E(n955), .CK(clk), .Q(\mem[17][5] ) );
  EDFFX1 \mem_reg[17][4]  ( .D(n894), .E(n955), .CK(clk), .Q(\mem[17][4] ) );
  EDFFX1 \mem_reg[17][3]  ( .D(n889), .E(n955), .CK(clk), .Q(\mem[17][3] ) );
  EDFFX1 \mem_reg[17][2]  ( .D(n884), .E(n955), .CK(clk), .Q(\mem[17][2] ) );
  EDFFX1 \mem_reg[17][1]  ( .D(n879), .E(n955), .CK(clk), .Q(\mem[17][1] ) );
  EDFFX1 \mem_reg[17][0]  ( .D(n874), .E(n955), .CK(clk), .Q(\mem[17][0] ) );
  EDFFX1 \mem_reg[21][7]  ( .D(data_in[7]), .E(n964), .CK(clk), .Q(
        \mem[21][7] ) );
  EDFFX1 \mem_reg[21][6]  ( .D(data_in[6]), .E(n964), .CK(clk), .Q(
        \mem[21][6] ) );
  EDFFX1 \mem_reg[21][5]  ( .D(data_in[5]), .E(n964), .CK(clk), .Q(
        \mem[21][5] ) );
  EDFFX1 \mem_reg[21][4]  ( .D(data_in[4]), .E(n964), .CK(clk), .Q(
        \mem[21][4] ) );
  EDFFX1 \mem_reg[21][3]  ( .D(data_in[3]), .E(n964), .CK(clk), .Q(
        \mem[21][3] ) );
  EDFFX1 \mem_reg[21][2]  ( .D(data_in[2]), .E(n964), .CK(clk), .Q(
        \mem[21][2] ) );
  EDFFX1 \mem_reg[21][1]  ( .D(data_in[1]), .E(n964), .CK(clk), .Q(
        \mem[21][1] ) );
  EDFFX1 \mem_reg[21][0]  ( .D(data_in[0]), .E(n964), .CK(clk), .Q(
        \mem[21][0] ) );
  EDFFX1 \mem_reg[25][7]  ( .D(data_in[7]), .E(n973), .CK(clk), .Q(
        \mem[25][7] ) );
  EDFFX1 \mem_reg[25][6]  ( .D(data_in[6]), .E(n973), .CK(clk), .Q(
        \mem[25][6] ) );
  EDFFX1 \mem_reg[25][5]  ( .D(data_in[5]), .E(n973), .CK(clk), .Q(
        \mem[25][5] ) );
  EDFFX1 \mem_reg[25][4]  ( .D(data_in[4]), .E(n973), .CK(clk), .Q(
        \mem[25][4] ) );
  EDFFX1 \mem_reg[25][3]  ( .D(data_in[3]), .E(n973), .CK(clk), .Q(
        \mem[25][3] ) );
  EDFFX1 \mem_reg[25][2]  ( .D(data_in[2]), .E(n973), .CK(clk), .Q(
        \mem[25][2] ) );
  EDFFX1 \mem_reg[25][1]  ( .D(data_in[1]), .E(n973), .CK(clk), .Q(
        \mem[25][1] ) );
  EDFFX1 \mem_reg[25][0]  ( .D(data_in[0]), .E(n973), .CK(clk), .Q(
        \mem[25][0] ) );
  EDFFX1 \mem_reg[29][7]  ( .D(data_in[7]), .E(n982), .CK(clk), .Q(
        \mem[29][7] ) );
  EDFFX1 \mem_reg[29][6]  ( .D(data_in[6]), .E(n982), .CK(clk), .Q(
        \mem[29][6] ) );
  EDFFX1 \mem_reg[29][5]  ( .D(data_in[5]), .E(n982), .CK(clk), .Q(
        \mem[29][5] ) );
  EDFFX1 \mem_reg[29][4]  ( .D(data_in[4]), .E(n982), .CK(clk), .Q(
        \mem[29][4] ) );
  EDFFX1 \mem_reg[29][3]  ( .D(data_in[3]), .E(n982), .CK(clk), .Q(
        \mem[29][3] ) );
  EDFFX1 \mem_reg[29][2]  ( .D(data_in[2]), .E(n982), .CK(clk), .Q(
        \mem[29][2] ) );
  EDFFX1 \mem_reg[29][1]  ( .D(data_in[1]), .E(n982), .CK(clk), .Q(
        \mem[29][1] ) );
  EDFFX1 \mem_reg[29][0]  ( .D(data_in[0]), .E(n982), .CK(clk), .Q(
        \mem[29][0] ) );
  EDFFX1 \mem_reg[33][7]  ( .D(n911), .E(n954), .CK(clk), .Q(\mem[33][7] ) );
  EDFFX1 \mem_reg[33][6]  ( .D(n906), .E(n954), .CK(clk), .Q(\mem[33][6] ) );
  EDFFX1 \mem_reg[33][5]  ( .D(n901), .E(n954), .CK(clk), .Q(\mem[33][5] ) );
  EDFFX1 \mem_reg[33][4]  ( .D(n896), .E(n954), .CK(clk), .Q(\mem[33][4] ) );
  EDFFX1 \mem_reg[33][3]  ( .D(n891), .E(n954), .CK(clk), .Q(\mem[33][3] ) );
  EDFFX1 \mem_reg[33][2]  ( .D(n886), .E(n954), .CK(clk), .Q(\mem[33][2] ) );
  EDFFX1 \mem_reg[33][1]  ( .D(n881), .E(n954), .CK(clk), .Q(\mem[33][1] ) );
  EDFFX1 \mem_reg[33][0]  ( .D(n876), .E(n954), .CK(clk), .Q(\mem[33][0] ) );
  EDFFX1 \mem_reg[37][7]  ( .D(n911), .E(n963), .CK(clk), .Q(\mem[37][7] ) );
  EDFFX1 \mem_reg[37][6]  ( .D(n906), .E(n963), .CK(clk), .Q(\mem[37][6] ) );
  EDFFX1 \mem_reg[37][5]  ( .D(n901), .E(n963), .CK(clk), .Q(\mem[37][5] ) );
  EDFFX1 \mem_reg[37][4]  ( .D(n896), .E(n963), .CK(clk), .Q(\mem[37][4] ) );
  EDFFX1 \mem_reg[37][3]  ( .D(n891), .E(n963), .CK(clk), .Q(\mem[37][3] ) );
  EDFFX1 \mem_reg[37][2]  ( .D(n886), .E(n963), .CK(clk), .Q(\mem[37][2] ) );
  EDFFX1 \mem_reg[37][1]  ( .D(n881), .E(n963), .CK(clk), .Q(\mem[37][1] ) );
  EDFFX1 \mem_reg[37][0]  ( .D(n876), .E(n963), .CK(clk), .Q(\mem[37][0] ) );
  EDFFX1 \mem_reg[41][7]  ( .D(n911), .E(n972), .CK(clk), .Q(\mem[41][7] ) );
  EDFFX1 \mem_reg[41][6]  ( .D(n906), .E(n972), .CK(clk), .Q(\mem[41][6] ) );
  EDFFX1 \mem_reg[41][5]  ( .D(n901), .E(n972), .CK(clk), .Q(\mem[41][5] ) );
  EDFFX1 \mem_reg[41][4]  ( .D(n896), .E(n972), .CK(clk), .Q(\mem[41][4] ) );
  EDFFX1 \mem_reg[41][3]  ( .D(n891), .E(n972), .CK(clk), .Q(\mem[41][3] ) );
  EDFFX1 \mem_reg[41][2]  ( .D(n886), .E(n972), .CK(clk), .Q(\mem[41][2] ) );
  EDFFX1 \mem_reg[41][1]  ( .D(n881), .E(n972), .CK(clk), .Q(\mem[41][1] ) );
  EDFFX1 \mem_reg[41][0]  ( .D(n876), .E(n972), .CK(clk), .Q(\mem[41][0] ) );
  EDFFX1 \mem_reg[45][7]  ( .D(n910), .E(n981), .CK(clk), .Q(\mem[45][7] ) );
  EDFFX1 \mem_reg[45][6]  ( .D(n905), .E(n981), .CK(clk), .Q(\mem[45][6] ) );
  EDFFX1 \mem_reg[45][5]  ( .D(n900), .E(n981), .CK(clk), .Q(\mem[45][5] ) );
  EDFFX1 \mem_reg[45][4]  ( .D(n895), .E(n981), .CK(clk), .Q(\mem[45][4] ) );
  EDFFX1 \mem_reg[45][3]  ( .D(n890), .E(n981), .CK(clk), .Q(\mem[45][3] ) );
  EDFFX1 \mem_reg[45][2]  ( .D(n885), .E(n981), .CK(clk), .Q(\mem[45][2] ) );
  EDFFX1 \mem_reg[45][1]  ( .D(n880), .E(n981), .CK(clk), .Q(\mem[45][1] ) );
  EDFFX1 \mem_reg[45][0]  ( .D(n875), .E(n981), .CK(clk), .Q(\mem[45][0] ) );
  EDFFX1 \mem_reg[49][7]  ( .D(n907), .E(n953), .CK(clk), .Q(\mem[49][7] ) );
  EDFFX1 \mem_reg[49][6]  ( .D(n902), .E(n953), .CK(clk), .Q(\mem[49][6] ) );
  EDFFX1 \mem_reg[49][5]  ( .D(n897), .E(n953), .CK(clk), .Q(\mem[49][5] ) );
  EDFFX1 \mem_reg[49][4]  ( .D(n892), .E(n953), .CK(clk), .Q(\mem[49][4] ) );
  EDFFX1 \mem_reg[49][3]  ( .D(n887), .E(n953), .CK(clk), .Q(\mem[49][3] ) );
  EDFFX1 \mem_reg[49][2]  ( .D(n882), .E(n953), .CK(clk), .Q(\mem[49][2] ) );
  EDFFX1 \mem_reg[49][1]  ( .D(n877), .E(n953), .CK(clk), .Q(\mem[49][1] ) );
  EDFFX1 \mem_reg[49][0]  ( .D(n872), .E(n953), .CK(clk), .Q(\mem[49][0] ) );
  EDFFX1 \mem_reg[53][7]  ( .D(n907), .E(n962), .CK(clk), .Q(\mem[53][7] ) );
  EDFFX1 \mem_reg[53][6]  ( .D(n902), .E(n962), .CK(clk), .Q(\mem[53][6] ) );
  EDFFX1 \mem_reg[53][5]  ( .D(n897), .E(n962), .CK(clk), .Q(\mem[53][5] ) );
  EDFFX1 \mem_reg[53][4]  ( .D(n892), .E(n962), .CK(clk), .Q(\mem[53][4] ) );
  EDFFX1 \mem_reg[53][3]  ( .D(n887), .E(n962), .CK(clk), .Q(\mem[53][3] ) );
  EDFFX1 \mem_reg[53][2]  ( .D(n882), .E(n962), .CK(clk), .Q(\mem[53][2] ) );
  EDFFX1 \mem_reg[53][1]  ( .D(n877), .E(n962), .CK(clk), .Q(\mem[53][1] ) );
  EDFFX1 \mem_reg[53][0]  ( .D(n872), .E(n962), .CK(clk), .Q(\mem[53][0] ) );
  EDFFX1 \mem_reg[57][7]  ( .D(n910), .E(n971), .CK(clk), .Q(\mem[57][7] ) );
  EDFFX1 \mem_reg[57][6]  ( .D(n905), .E(n971), .CK(clk), .Q(\mem[57][6] ) );
  EDFFX1 \mem_reg[57][5]  ( .D(n900), .E(n971), .CK(clk), .Q(\mem[57][5] ) );
  EDFFX1 \mem_reg[57][4]  ( .D(n895), .E(n971), .CK(clk), .Q(\mem[57][4] ) );
  EDFFX1 \mem_reg[57][3]  ( .D(n890), .E(n971), .CK(clk), .Q(\mem[57][3] ) );
  EDFFX1 \mem_reg[57][2]  ( .D(n885), .E(n971), .CK(clk), .Q(\mem[57][2] ) );
  EDFFX1 \mem_reg[57][1]  ( .D(n880), .E(n971), .CK(clk), .Q(\mem[57][1] ) );
  EDFFX1 \mem_reg[57][0]  ( .D(n875), .E(n971), .CK(clk), .Q(\mem[57][0] ) );
  EDFFX1 \mem_reg[61][7]  ( .D(n910), .E(n980), .CK(clk), .Q(\mem[61][7] ) );
  EDFFX1 \mem_reg[61][6]  ( .D(n905), .E(n980), .CK(clk), .Q(\mem[61][6] ) );
  EDFFX1 \mem_reg[61][5]  ( .D(n900), .E(n980), .CK(clk), .Q(\mem[61][5] ) );
  EDFFX1 \mem_reg[61][4]  ( .D(n895), .E(n980), .CK(clk), .Q(\mem[61][4] ) );
  EDFFX1 \mem_reg[61][3]  ( .D(n890), .E(n980), .CK(clk), .Q(\mem[61][3] ) );
  EDFFX1 \mem_reg[61][2]  ( .D(n885), .E(n980), .CK(clk), .Q(\mem[61][2] ) );
  EDFFX1 \mem_reg[61][1]  ( .D(n880), .E(n980), .CK(clk), .Q(\mem[61][1] ) );
  EDFFX1 \mem_reg[61][0]  ( .D(n875), .E(n980), .CK(clk), .Q(\mem[61][0] ) );
  EDFFX1 \mem_reg[65][7]  ( .D(n910), .E(n952), .CK(clk), .Q(\mem[65][7] ) );
  EDFFX1 \mem_reg[65][6]  ( .D(n905), .E(n952), .CK(clk), .Q(\mem[65][6] ) );
  EDFFX1 \mem_reg[65][5]  ( .D(n900), .E(n952), .CK(clk), .Q(\mem[65][5] ) );
  EDFFX1 \mem_reg[65][4]  ( .D(n895), .E(n952), .CK(clk), .Q(\mem[65][4] ) );
  EDFFX1 \mem_reg[65][3]  ( .D(n890), .E(n952), .CK(clk), .Q(\mem[65][3] ) );
  EDFFX1 \mem_reg[65][2]  ( .D(n885), .E(n952), .CK(clk), .Q(\mem[65][2] ) );
  EDFFX1 \mem_reg[65][1]  ( .D(n880), .E(n952), .CK(clk), .Q(\mem[65][1] ) );
  EDFFX1 \mem_reg[65][0]  ( .D(n875), .E(n952), .CK(clk), .Q(\mem[65][0] ) );
  EDFFX1 \mem_reg[69][7]  ( .D(n907), .E(n961), .CK(clk), .Q(\mem[69][7] ) );
  EDFFX1 \mem_reg[69][6]  ( .D(n902), .E(n961), .CK(clk), .Q(\mem[69][6] ) );
  EDFFX1 \mem_reg[69][5]  ( .D(n897), .E(n961), .CK(clk), .Q(\mem[69][5] ) );
  EDFFX1 \mem_reg[69][4]  ( .D(n892), .E(n961), .CK(clk), .Q(\mem[69][4] ) );
  EDFFX1 \mem_reg[69][3]  ( .D(n887), .E(n961), .CK(clk), .Q(\mem[69][3] ) );
  EDFFX1 \mem_reg[69][2]  ( .D(n882), .E(n961), .CK(clk), .Q(\mem[69][2] ) );
  EDFFX1 \mem_reg[69][1]  ( .D(n877), .E(n961), .CK(clk), .Q(\mem[69][1] ) );
  EDFFX1 \mem_reg[69][0]  ( .D(n872), .E(n961), .CK(clk), .Q(\mem[69][0] ) );
  EDFFX1 \mem_reg[73][7]  ( .D(n909), .E(n970), .CK(clk), .Q(\mem[73][7] ) );
  EDFFX1 \mem_reg[73][6]  ( .D(n904), .E(n970), .CK(clk), .Q(\mem[73][6] ) );
  EDFFX1 \mem_reg[73][5]  ( .D(n899), .E(n970), .CK(clk), .Q(\mem[73][5] ) );
  EDFFX1 \mem_reg[73][4]  ( .D(n894), .E(n970), .CK(clk), .Q(\mem[73][4] ) );
  EDFFX1 \mem_reg[73][3]  ( .D(n889), .E(n970), .CK(clk), .Q(\mem[73][3] ) );
  EDFFX1 \mem_reg[73][2]  ( .D(n884), .E(n970), .CK(clk), .Q(\mem[73][2] ) );
  EDFFX1 \mem_reg[73][1]  ( .D(n879), .E(n970), .CK(clk), .Q(\mem[73][1] ) );
  EDFFX1 \mem_reg[73][0]  ( .D(n874), .E(n970), .CK(clk), .Q(\mem[73][0] ) );
  EDFFX1 \mem_reg[77][7]  ( .D(n910), .E(n979), .CK(clk), .Q(\mem[77][7] ) );
  EDFFX1 \mem_reg[77][6]  ( .D(n905), .E(n979), .CK(clk), .Q(\mem[77][6] ) );
  EDFFX1 \mem_reg[77][5]  ( .D(n900), .E(n979), .CK(clk), .Q(\mem[77][5] ) );
  EDFFX1 \mem_reg[77][4]  ( .D(n895), .E(n979), .CK(clk), .Q(\mem[77][4] ) );
  EDFFX1 \mem_reg[77][3]  ( .D(n890), .E(n979), .CK(clk), .Q(\mem[77][3] ) );
  EDFFX1 \mem_reg[77][2]  ( .D(n885), .E(n979), .CK(clk), .Q(\mem[77][2] ) );
  EDFFX1 \mem_reg[77][1]  ( .D(n880), .E(n979), .CK(clk), .Q(\mem[77][1] ) );
  EDFFX1 \mem_reg[77][0]  ( .D(n875), .E(n979), .CK(clk), .Q(\mem[77][0] ) );
  EDFFX1 \mem_reg[81][7]  ( .D(n909), .E(n951), .CK(clk), .Q(\mem[81][7] ) );
  EDFFX1 \mem_reg[81][6]  ( .D(n904), .E(n951), .CK(clk), .Q(\mem[81][6] ) );
  EDFFX1 \mem_reg[81][5]  ( .D(n899), .E(n951), .CK(clk), .Q(\mem[81][5] ) );
  EDFFX1 \mem_reg[81][4]  ( .D(n894), .E(n951), .CK(clk), .Q(\mem[81][4] ) );
  EDFFX1 \mem_reg[81][3]  ( .D(n889), .E(n951), .CK(clk), .Q(\mem[81][3] ) );
  EDFFX1 \mem_reg[81][2]  ( .D(n884), .E(n951), .CK(clk), .Q(\mem[81][2] ) );
  EDFFX1 \mem_reg[81][1]  ( .D(n879), .E(n951), .CK(clk), .Q(\mem[81][1] ) );
  EDFFX1 \mem_reg[81][0]  ( .D(n874), .E(n951), .CK(clk), .Q(\mem[81][0] ) );
  EDFFX1 \mem_reg[85][7]  ( .D(n909), .E(n960), .CK(clk), .Q(\mem[85][7] ) );
  EDFFX1 \mem_reg[85][6]  ( .D(n904), .E(n960), .CK(clk), .Q(\mem[85][6] ) );
  EDFFX1 \mem_reg[85][5]  ( .D(n899), .E(n960), .CK(clk), .Q(\mem[85][5] ) );
  EDFFX1 \mem_reg[85][4]  ( .D(n894), .E(n960), .CK(clk), .Q(\mem[85][4] ) );
  EDFFX1 \mem_reg[85][3]  ( .D(n889), .E(n960), .CK(clk), .Q(\mem[85][3] ) );
  EDFFX1 \mem_reg[85][2]  ( .D(n884), .E(n960), .CK(clk), .Q(\mem[85][2] ) );
  EDFFX1 \mem_reg[85][1]  ( .D(n879), .E(n960), .CK(clk), .Q(\mem[85][1] ) );
  EDFFX1 \mem_reg[85][0]  ( .D(n874), .E(n960), .CK(clk), .Q(\mem[85][0] ) );
  EDFFX1 \mem_reg[89][7]  ( .D(n909), .E(n969), .CK(clk), .Q(\mem[89][7] ) );
  EDFFX1 \mem_reg[89][6]  ( .D(n904), .E(n969), .CK(clk), .Q(\mem[89][6] ) );
  EDFFX1 \mem_reg[89][5]  ( .D(n899), .E(n969), .CK(clk), .Q(\mem[89][5] ) );
  EDFFX1 \mem_reg[89][4]  ( .D(n894), .E(n969), .CK(clk), .Q(\mem[89][4] ) );
  EDFFX1 \mem_reg[89][3]  ( .D(n889), .E(n969), .CK(clk), .Q(\mem[89][3] ) );
  EDFFX1 \mem_reg[89][2]  ( .D(n884), .E(n969), .CK(clk), .Q(\mem[89][2] ) );
  EDFFX1 \mem_reg[89][1]  ( .D(n879), .E(n969), .CK(clk), .Q(\mem[89][1] ) );
  EDFFX1 \mem_reg[89][0]  ( .D(n874), .E(n969), .CK(clk), .Q(\mem[89][0] ) );
  EDFFX1 \mem_reg[93][7]  ( .D(n908), .E(n978), .CK(clk), .Q(\mem[93][7] ) );
  EDFFX1 \mem_reg[93][6]  ( .D(n903), .E(n978), .CK(clk), .Q(\mem[93][6] ) );
  EDFFX1 \mem_reg[93][5]  ( .D(n898), .E(n978), .CK(clk), .Q(\mem[93][5] ) );
  EDFFX1 \mem_reg[93][4]  ( .D(n893), .E(n978), .CK(clk), .Q(\mem[93][4] ) );
  EDFFX1 \mem_reg[93][3]  ( .D(n888), .E(n978), .CK(clk), .Q(\mem[93][3] ) );
  EDFFX1 \mem_reg[93][2]  ( .D(n883), .E(n978), .CK(clk), .Q(\mem[93][2] ) );
  EDFFX1 \mem_reg[93][1]  ( .D(n878), .E(n978), .CK(clk), .Q(\mem[93][1] ) );
  EDFFX1 \mem_reg[93][0]  ( .D(n873), .E(n978), .CK(clk), .Q(\mem[93][0] ) );
  EDFFX1 \mem_reg[97][7]  ( .D(n911), .E(n950), .CK(clk), .Q(\mem[97][7] ) );
  EDFFX1 \mem_reg[97][6]  ( .D(n906), .E(n950), .CK(clk), .Q(\mem[97][6] ) );
  EDFFX1 \mem_reg[97][5]  ( .D(n901), .E(n950), .CK(clk), .Q(\mem[97][5] ) );
  EDFFX1 \mem_reg[97][4]  ( .D(n896), .E(n950), .CK(clk), .Q(\mem[97][4] ) );
  EDFFX1 \mem_reg[97][3]  ( .D(n891), .E(n950), .CK(clk), .Q(\mem[97][3] ) );
  EDFFX1 \mem_reg[97][2]  ( .D(n886), .E(n950), .CK(clk), .Q(\mem[97][2] ) );
  EDFFX1 \mem_reg[97][1]  ( .D(n881), .E(n950), .CK(clk), .Q(\mem[97][1] ) );
  EDFFX1 \mem_reg[97][0]  ( .D(n876), .E(n950), .CK(clk), .Q(\mem[97][0] ) );
  EDFFX1 \mem_reg[101][7]  ( .D(n910), .E(n959), .CK(clk), .Q(\mem[101][7] )
         );
  EDFFX1 \mem_reg[101][6]  ( .D(n905), .E(n959), .CK(clk), .Q(\mem[101][6] )
         );
  EDFFX1 \mem_reg[101][5]  ( .D(n900), .E(n959), .CK(clk), .Q(\mem[101][5] )
         );
  EDFFX1 \mem_reg[101][4]  ( .D(n895), .E(n959), .CK(clk), .Q(\mem[101][4] )
         );
  EDFFX1 \mem_reg[101][3]  ( .D(n890), .E(n959), .CK(clk), .Q(\mem[101][3] )
         );
  EDFFX1 \mem_reg[101][2]  ( .D(n885), .E(n959), .CK(clk), .Q(\mem[101][2] )
         );
  EDFFX1 \mem_reg[101][1]  ( .D(n880), .E(n959), .CK(clk), .Q(\mem[101][1] )
         );
  EDFFX1 \mem_reg[101][0]  ( .D(n875), .E(n959), .CK(clk), .Q(\mem[101][0] )
         );
  EDFFX1 \mem_reg[105][7]  ( .D(n908), .E(n968), .CK(clk), .Q(\mem[105][7] )
         );
  EDFFX1 \mem_reg[105][6]  ( .D(n903), .E(n968), .CK(clk), .Q(\mem[105][6] )
         );
  EDFFX1 \mem_reg[105][5]  ( .D(n898), .E(n968), .CK(clk), .Q(\mem[105][5] )
         );
  EDFFX1 \mem_reg[105][4]  ( .D(n893), .E(n968), .CK(clk), .Q(\mem[105][4] )
         );
  EDFFX1 \mem_reg[105][3]  ( .D(n888), .E(n968), .CK(clk), .Q(\mem[105][3] )
         );
  EDFFX1 \mem_reg[105][2]  ( .D(n883), .E(n968), .CK(clk), .Q(\mem[105][2] )
         );
  EDFFX1 \mem_reg[105][1]  ( .D(n878), .E(n968), .CK(clk), .Q(\mem[105][1] )
         );
  EDFFX1 \mem_reg[105][0]  ( .D(n873), .E(n968), .CK(clk), .Q(\mem[105][0] )
         );
  EDFFX1 \mem_reg[109][7]  ( .D(n908), .E(n977), .CK(clk), .Q(\mem[109][7] )
         );
  EDFFX1 \mem_reg[109][6]  ( .D(n903), .E(n977), .CK(clk), .Q(\mem[109][6] )
         );
  EDFFX1 \mem_reg[109][5]  ( .D(n898), .E(n977), .CK(clk), .Q(\mem[109][5] )
         );
  EDFFX1 \mem_reg[109][4]  ( .D(n893), .E(n977), .CK(clk), .Q(\mem[109][4] )
         );
  EDFFX1 \mem_reg[109][3]  ( .D(n888), .E(n977), .CK(clk), .Q(\mem[109][3] )
         );
  EDFFX1 \mem_reg[109][2]  ( .D(n883), .E(n977), .CK(clk), .Q(\mem[109][2] )
         );
  EDFFX1 \mem_reg[109][1]  ( .D(n878), .E(n977), .CK(clk), .Q(\mem[109][1] )
         );
  EDFFX1 \mem_reg[109][0]  ( .D(n873), .E(n977), .CK(clk), .Q(\mem[109][0] )
         );
  EDFFX1 \mem_reg[113][7]  ( .D(n908), .E(n949), .CK(clk), .Q(\mem[113][7] )
         );
  EDFFX1 \mem_reg[113][6]  ( .D(n903), .E(n949), .CK(clk), .Q(\mem[113][6] )
         );
  EDFFX1 \mem_reg[113][5]  ( .D(n898), .E(n949), .CK(clk), .Q(\mem[113][5] )
         );
  EDFFX1 \mem_reg[113][4]  ( .D(n893), .E(n949), .CK(clk), .Q(\mem[113][4] )
         );
  EDFFX1 \mem_reg[113][3]  ( .D(n888), .E(n949), .CK(clk), .Q(\mem[113][3] )
         );
  EDFFX1 \mem_reg[113][2]  ( .D(n883), .E(n949), .CK(clk), .Q(\mem[113][2] )
         );
  EDFFX1 \mem_reg[113][1]  ( .D(n878), .E(n949), .CK(clk), .Q(\mem[113][1] )
         );
  EDFFX1 \mem_reg[113][0]  ( .D(n873), .E(n949), .CK(clk), .Q(\mem[113][0] )
         );
  EDFFX1 \mem_reg[117][7]  ( .D(n907), .E(n958), .CK(clk), .Q(\mem[117][7] )
         );
  EDFFX1 \mem_reg[117][6]  ( .D(n902), .E(n958), .CK(clk), .Q(\mem[117][6] )
         );
  EDFFX1 \mem_reg[117][5]  ( .D(n897), .E(n958), .CK(clk), .Q(\mem[117][5] )
         );
  EDFFX1 \mem_reg[117][4]  ( .D(n892), .E(n958), .CK(clk), .Q(\mem[117][4] )
         );
  EDFFX1 \mem_reg[117][3]  ( .D(n887), .E(n958), .CK(clk), .Q(\mem[117][3] )
         );
  EDFFX1 \mem_reg[117][2]  ( .D(n882), .E(n958), .CK(clk), .Q(\mem[117][2] )
         );
  EDFFX1 \mem_reg[117][1]  ( .D(n877), .E(n958), .CK(clk), .Q(\mem[117][1] )
         );
  EDFFX1 \mem_reg[117][0]  ( .D(n872), .E(n958), .CK(clk), .Q(\mem[117][0] )
         );
  EDFFX1 \mem_reg[121][7]  ( .D(n907), .E(n967), .CK(clk), .Q(\mem[121][7] )
         );
  EDFFX1 \mem_reg[121][6]  ( .D(n902), .E(n967), .CK(clk), .Q(\mem[121][6] )
         );
  EDFFX1 \mem_reg[121][5]  ( .D(n897), .E(n967), .CK(clk), .Q(\mem[121][5] )
         );
  EDFFX1 \mem_reg[121][4]  ( .D(n892), .E(n967), .CK(clk), .Q(\mem[121][4] )
         );
  EDFFX1 \mem_reg[121][3]  ( .D(n887), .E(n967), .CK(clk), .Q(\mem[121][3] )
         );
  EDFFX1 \mem_reg[121][2]  ( .D(n882), .E(n967), .CK(clk), .Q(\mem[121][2] )
         );
  EDFFX1 \mem_reg[121][1]  ( .D(n877), .E(n967), .CK(clk), .Q(\mem[121][1] )
         );
  EDFFX1 \mem_reg[121][0]  ( .D(n872), .E(n967), .CK(clk), .Q(\mem[121][0] )
         );
  EDFFX1 \mem_reg[125][7]  ( .D(n907), .E(n976), .CK(clk), .Q(\mem[125][7] )
         );
  EDFFX1 \mem_reg[125][6]  ( .D(n902), .E(n976), .CK(clk), .Q(\mem[125][6] )
         );
  EDFFX1 \mem_reg[125][5]  ( .D(n897), .E(n976), .CK(clk), .Q(\mem[125][5] )
         );
  EDFFX1 \mem_reg[125][4]  ( .D(n892), .E(n976), .CK(clk), .Q(\mem[125][4] )
         );
  EDFFX1 \mem_reg[125][3]  ( .D(n887), .E(n976), .CK(clk), .Q(\mem[125][3] )
         );
  EDFFX1 \mem_reg[125][2]  ( .D(n882), .E(n976), .CK(clk), .Q(\mem[125][2] )
         );
  EDFFX1 \mem_reg[125][1]  ( .D(n877), .E(n976), .CK(clk), .Q(\mem[125][1] )
         );
  EDFFX1 \mem_reg[125][0]  ( .D(n872), .E(n976), .CK(clk), .Q(\mem[125][0] )
         );
  EDFFX1 \mem_reg[3][7]  ( .D(n910), .E(n920), .CK(clk), .Q(\mem[3][7] ) );
  EDFFX1 \mem_reg[3][6]  ( .D(n905), .E(n920), .CK(clk), .Q(\mem[3][6] ) );
  EDFFX1 \mem_reg[3][5]  ( .D(n900), .E(n920), .CK(clk), .Q(\mem[3][5] ) );
  EDFFX1 \mem_reg[3][4]  ( .D(n895), .E(n920), .CK(clk), .Q(\mem[3][4] ) );
  EDFFX1 \mem_reg[3][3]  ( .D(n890), .E(n920), .CK(clk), .Q(\mem[3][3] ) );
  EDFFX1 \mem_reg[3][2]  ( .D(n885), .E(n920), .CK(clk), .Q(\mem[3][2] ) );
  EDFFX1 \mem_reg[3][1]  ( .D(n880), .E(n920), .CK(clk), .Q(\mem[3][1] ) );
  EDFFX1 \mem_reg[3][0]  ( .D(n875), .E(n920), .CK(clk), .Q(\mem[3][0] ) );
  EDFFX1 \mem_reg[7][7]  ( .D(n907), .E(n929), .CK(clk), .Q(\mem[7][7] ) );
  EDFFX1 \mem_reg[7][6]  ( .D(n902), .E(n929), .CK(clk), .Q(\mem[7][6] ) );
  EDFFX1 \mem_reg[7][5]  ( .D(n897), .E(n929), .CK(clk), .Q(\mem[7][5] ) );
  EDFFX1 \mem_reg[7][4]  ( .D(n892), .E(n929), .CK(clk), .Q(\mem[7][4] ) );
  EDFFX1 \mem_reg[7][3]  ( .D(n887), .E(n929), .CK(clk), .Q(\mem[7][3] ) );
  EDFFX1 \mem_reg[7][2]  ( .D(n882), .E(n929), .CK(clk), .Q(\mem[7][2] ) );
  EDFFX1 \mem_reg[7][1]  ( .D(n877), .E(n929), .CK(clk), .Q(\mem[7][1] ) );
  EDFFX1 \mem_reg[7][0]  ( .D(n872), .E(n929), .CK(clk), .Q(\mem[7][0] ) );
  EDFFX1 \mem_reg[11][7]  ( .D(n910), .E(n938), .CK(clk), .Q(\mem[11][7] ) );
  EDFFX1 \mem_reg[11][6]  ( .D(n905), .E(n938), .CK(clk), .Q(\mem[11][6] ) );
  EDFFX1 \mem_reg[11][5]  ( .D(n900), .E(n938), .CK(clk), .Q(\mem[11][5] ) );
  EDFFX1 \mem_reg[11][4]  ( .D(n895), .E(n938), .CK(clk), .Q(\mem[11][4] ) );
  EDFFX1 \mem_reg[11][3]  ( .D(n890), .E(n938), .CK(clk), .Q(\mem[11][3] ) );
  EDFFX1 \mem_reg[11][2]  ( .D(n885), .E(n938), .CK(clk), .Q(\mem[11][2] ) );
  EDFFX1 \mem_reg[11][1]  ( .D(n880), .E(n938), .CK(clk), .Q(\mem[11][1] ) );
  EDFFX1 \mem_reg[11][0]  ( .D(n875), .E(n938), .CK(clk), .Q(\mem[11][0] ) );
  EDFFX1 \mem_reg[15][7]  ( .D(n909), .E(n947), .CK(clk), .Q(\mem[15][7] ) );
  EDFFX1 \mem_reg[15][6]  ( .D(n904), .E(n947), .CK(clk), .Q(\mem[15][6] ) );
  EDFFX1 \mem_reg[15][5]  ( .D(n899), .E(n947), .CK(clk), .Q(\mem[15][5] ) );
  EDFFX1 \mem_reg[15][4]  ( .D(n894), .E(n947), .CK(clk), .Q(\mem[15][4] ) );
  EDFFX1 \mem_reg[15][3]  ( .D(n889), .E(n947), .CK(clk), .Q(\mem[15][3] ) );
  EDFFX1 \mem_reg[15][2]  ( .D(n884), .E(n947), .CK(clk), .Q(\mem[15][2] ) );
  EDFFX1 \mem_reg[15][1]  ( .D(n879), .E(n947), .CK(clk), .Q(\mem[15][1] ) );
  EDFFX1 \mem_reg[15][0]  ( .D(n874), .E(n947), .CK(clk), .Q(\mem[15][0] ) );
  EDFFX1 \mem_reg[19][7]  ( .D(data_in[7]), .E(n919), .CK(clk), .Q(
        \mem[19][7] ) );
  EDFFX1 \mem_reg[19][6]  ( .D(data_in[6]), .E(n919), .CK(clk), .Q(
        \mem[19][6] ) );
  EDFFX1 \mem_reg[19][5]  ( .D(data_in[5]), .E(n919), .CK(clk), .Q(
        \mem[19][5] ) );
  EDFFX1 \mem_reg[19][4]  ( .D(data_in[4]), .E(n919), .CK(clk), .Q(
        \mem[19][4] ) );
  EDFFX1 \mem_reg[19][3]  ( .D(data_in[3]), .E(n919), .CK(clk), .Q(
        \mem[19][3] ) );
  EDFFX1 \mem_reg[19][2]  ( .D(data_in[2]), .E(n919), .CK(clk), .Q(
        \mem[19][2] ) );
  EDFFX1 \mem_reg[19][1]  ( .D(data_in[1]), .E(n919), .CK(clk), .Q(
        \mem[19][1] ) );
  EDFFX1 \mem_reg[19][0]  ( .D(data_in[0]), .E(n919), .CK(clk), .Q(
        \mem[19][0] ) );
  EDFFX1 \mem_reg[23][7]  ( .D(data_in[7]), .E(n928), .CK(clk), .Q(
        \mem[23][7] ) );
  EDFFX1 \mem_reg[23][6]  ( .D(data_in[6]), .E(n928), .CK(clk), .Q(
        \mem[23][6] ) );
  EDFFX1 \mem_reg[23][5]  ( .D(data_in[5]), .E(n928), .CK(clk), .Q(
        \mem[23][5] ) );
  EDFFX1 \mem_reg[23][4]  ( .D(data_in[4]), .E(n928), .CK(clk), .Q(
        \mem[23][4] ) );
  EDFFX1 \mem_reg[23][3]  ( .D(data_in[3]), .E(n928), .CK(clk), .Q(
        \mem[23][3] ) );
  EDFFX1 \mem_reg[23][2]  ( .D(data_in[2]), .E(n928), .CK(clk), .Q(
        \mem[23][2] ) );
  EDFFX1 \mem_reg[23][1]  ( .D(data_in[1]), .E(n928), .CK(clk), .Q(
        \mem[23][1] ) );
  EDFFX1 \mem_reg[23][0]  ( .D(data_in[0]), .E(n928), .CK(clk), .Q(
        \mem[23][0] ) );
  EDFFX1 \mem_reg[27][7]  ( .D(data_in[7]), .E(n937), .CK(clk), .Q(
        \mem[27][7] ) );
  EDFFX1 \mem_reg[27][6]  ( .D(data_in[6]), .E(n937), .CK(clk), .Q(
        \mem[27][6] ) );
  EDFFX1 \mem_reg[27][5]  ( .D(data_in[5]), .E(n937), .CK(clk), .Q(
        \mem[27][5] ) );
  EDFFX1 \mem_reg[27][4]  ( .D(data_in[4]), .E(n937), .CK(clk), .Q(
        \mem[27][4] ) );
  EDFFX1 \mem_reg[27][3]  ( .D(data_in[3]), .E(n937), .CK(clk), .Q(
        \mem[27][3] ) );
  EDFFX1 \mem_reg[27][2]  ( .D(data_in[2]), .E(n937), .CK(clk), .Q(
        \mem[27][2] ) );
  EDFFX1 \mem_reg[27][1]  ( .D(data_in[1]), .E(n937), .CK(clk), .Q(
        \mem[27][1] ) );
  EDFFX1 \mem_reg[27][0]  ( .D(data_in[0]), .E(n937), .CK(clk), .Q(
        \mem[27][0] ) );
  EDFFX1 \mem_reg[31][7]  ( .D(data_in[7]), .E(n946), .CK(clk), .Q(
        \mem[31][7] ) );
  EDFFX1 \mem_reg[31][6]  ( .D(data_in[6]), .E(n946), .CK(clk), .Q(
        \mem[31][6] ) );
  EDFFX1 \mem_reg[31][5]  ( .D(data_in[5]), .E(n946), .CK(clk), .Q(
        \mem[31][5] ) );
  EDFFX1 \mem_reg[31][4]  ( .D(data_in[4]), .E(n946), .CK(clk), .Q(
        \mem[31][4] ) );
  EDFFX1 \mem_reg[31][3]  ( .D(data_in[3]), .E(n946), .CK(clk), .Q(
        \mem[31][3] ) );
  EDFFX1 \mem_reg[31][2]  ( .D(data_in[2]), .E(n946), .CK(clk), .Q(
        \mem[31][2] ) );
  EDFFX1 \mem_reg[31][1]  ( .D(data_in[1]), .E(n946), .CK(clk), .Q(
        \mem[31][1] ) );
  EDFFX1 \mem_reg[31][0]  ( .D(data_in[0]), .E(n946), .CK(clk), .Q(
        \mem[31][0] ) );
  EDFFX1 \mem_reg[35][7]  ( .D(n911), .E(n918), .CK(clk), .Q(\mem[35][7] ) );
  EDFFX1 \mem_reg[35][6]  ( .D(n906), .E(n918), .CK(clk), .Q(\mem[35][6] ) );
  EDFFX1 \mem_reg[35][5]  ( .D(n901), .E(n918), .CK(clk), .Q(\mem[35][5] ) );
  EDFFX1 \mem_reg[35][4]  ( .D(n896), .E(n918), .CK(clk), .Q(\mem[35][4] ) );
  EDFFX1 \mem_reg[35][3]  ( .D(n891), .E(n918), .CK(clk), .Q(\mem[35][3] ) );
  EDFFX1 \mem_reg[35][2]  ( .D(n886), .E(n918), .CK(clk), .Q(\mem[35][2] ) );
  EDFFX1 \mem_reg[35][1]  ( .D(n881), .E(n918), .CK(clk), .Q(\mem[35][1] ) );
  EDFFX1 \mem_reg[35][0]  ( .D(n876), .E(n918), .CK(clk), .Q(\mem[35][0] ) );
  EDFFX1 \mem_reg[39][7]  ( .D(n911), .E(n927), .CK(clk), .Q(\mem[39][7] ) );
  EDFFX1 \mem_reg[39][6]  ( .D(n906), .E(n927), .CK(clk), .Q(\mem[39][6] ) );
  EDFFX1 \mem_reg[39][5]  ( .D(n901), .E(n927), .CK(clk), .Q(\mem[39][5] ) );
  EDFFX1 \mem_reg[39][4]  ( .D(n896), .E(n927), .CK(clk), .Q(\mem[39][4] ) );
  EDFFX1 \mem_reg[39][3]  ( .D(n891), .E(n927), .CK(clk), .Q(\mem[39][3] ) );
  EDFFX1 \mem_reg[39][2]  ( .D(n886), .E(n927), .CK(clk), .Q(\mem[39][2] ) );
  EDFFX1 \mem_reg[39][1]  ( .D(n881), .E(n927), .CK(clk), .Q(\mem[39][1] ) );
  EDFFX1 \mem_reg[39][0]  ( .D(n876), .E(n927), .CK(clk), .Q(\mem[39][0] ) );
  EDFFX1 \mem_reg[43][7]  ( .D(n911), .E(n936), .CK(clk), .Q(\mem[43][7] ) );
  EDFFX1 \mem_reg[43][6]  ( .D(n906), .E(n936), .CK(clk), .Q(\mem[43][6] ) );
  EDFFX1 \mem_reg[43][5]  ( .D(n901), .E(n936), .CK(clk), .Q(\mem[43][5] ) );
  EDFFX1 \mem_reg[43][4]  ( .D(n896), .E(n936), .CK(clk), .Q(\mem[43][4] ) );
  EDFFX1 \mem_reg[43][3]  ( .D(n891), .E(n936), .CK(clk), .Q(\mem[43][3] ) );
  EDFFX1 \mem_reg[43][2]  ( .D(n886), .E(n936), .CK(clk), .Q(\mem[43][2] ) );
  EDFFX1 \mem_reg[43][1]  ( .D(n881), .E(n936), .CK(clk), .Q(\mem[43][1] ) );
  EDFFX1 \mem_reg[43][0]  ( .D(n876), .E(n936), .CK(clk), .Q(\mem[43][0] ) );
  EDFFX1 \mem_reg[47][7]  ( .D(n908), .E(n945), .CK(clk), .Q(\mem[47][7] ) );
  EDFFX1 \mem_reg[47][6]  ( .D(n903), .E(n945), .CK(clk), .Q(\mem[47][6] ) );
  EDFFX1 \mem_reg[47][5]  ( .D(n898), .E(n945), .CK(clk), .Q(\mem[47][5] ) );
  EDFFX1 \mem_reg[47][4]  ( .D(n893), .E(n945), .CK(clk), .Q(\mem[47][4] ) );
  EDFFX1 \mem_reg[47][3]  ( .D(n888), .E(n945), .CK(clk), .Q(\mem[47][3] ) );
  EDFFX1 \mem_reg[47][2]  ( .D(n883), .E(n945), .CK(clk), .Q(\mem[47][2] ) );
  EDFFX1 \mem_reg[47][1]  ( .D(n878), .E(n945), .CK(clk), .Q(\mem[47][1] ) );
  EDFFX1 \mem_reg[47][0]  ( .D(n873), .E(n945), .CK(clk), .Q(\mem[47][0] ) );
  EDFFX1 \mem_reg[51][7]  ( .D(n907), .E(n917), .CK(clk), .Q(\mem[51][7] ) );
  EDFFX1 \mem_reg[51][6]  ( .D(n902), .E(n917), .CK(clk), .Q(\mem[51][6] ) );
  EDFFX1 \mem_reg[51][5]  ( .D(n897), .E(n917), .CK(clk), .Q(\mem[51][5] ) );
  EDFFX1 \mem_reg[51][4]  ( .D(n892), .E(n917), .CK(clk), .Q(\mem[51][4] ) );
  EDFFX1 \mem_reg[51][3]  ( .D(n887), .E(n917), .CK(clk), .Q(\mem[51][3] ) );
  EDFFX1 \mem_reg[51][2]  ( .D(n882), .E(n917), .CK(clk), .Q(\mem[51][2] ) );
  EDFFX1 \mem_reg[51][1]  ( .D(n877), .E(n917), .CK(clk), .Q(\mem[51][1] ) );
  EDFFX1 \mem_reg[51][0]  ( .D(n872), .E(n917), .CK(clk), .Q(\mem[51][0] ) );
  EDFFX1 \mem_reg[55][7]  ( .D(n911), .E(n926), .CK(clk), .Q(\mem[55][7] ) );
  EDFFX1 \mem_reg[55][6]  ( .D(n906), .E(n926), .CK(clk), .Q(\mem[55][6] ) );
  EDFFX1 \mem_reg[55][5]  ( .D(n901), .E(n926), .CK(clk), .Q(\mem[55][5] ) );
  EDFFX1 \mem_reg[55][4]  ( .D(n896), .E(n926), .CK(clk), .Q(\mem[55][4] ) );
  EDFFX1 \mem_reg[55][3]  ( .D(n891), .E(n926), .CK(clk), .Q(\mem[55][3] ) );
  EDFFX1 \mem_reg[55][2]  ( .D(n886), .E(n926), .CK(clk), .Q(\mem[55][2] ) );
  EDFFX1 \mem_reg[55][1]  ( .D(n881), .E(n926), .CK(clk), .Q(\mem[55][1] ) );
  EDFFX1 \mem_reg[55][0]  ( .D(n876), .E(n926), .CK(clk), .Q(\mem[55][0] ) );
  EDFFX1 \mem_reg[59][7]  ( .D(n910), .E(n935), .CK(clk), .Q(\mem[59][7] ) );
  EDFFX1 \mem_reg[59][6]  ( .D(n905), .E(n935), .CK(clk), .Q(\mem[59][6] ) );
  EDFFX1 \mem_reg[59][5]  ( .D(n900), .E(n935), .CK(clk), .Q(\mem[59][5] ) );
  EDFFX1 \mem_reg[59][4]  ( .D(n895), .E(n935), .CK(clk), .Q(\mem[59][4] ) );
  EDFFX1 \mem_reg[59][3]  ( .D(n890), .E(n935), .CK(clk), .Q(\mem[59][3] ) );
  EDFFX1 \mem_reg[59][2]  ( .D(n885), .E(n935), .CK(clk), .Q(\mem[59][2] ) );
  EDFFX1 \mem_reg[59][1]  ( .D(n880), .E(n935), .CK(clk), .Q(\mem[59][1] ) );
  EDFFX1 \mem_reg[59][0]  ( .D(n875), .E(n935), .CK(clk), .Q(\mem[59][0] ) );
  EDFFX1 \mem_reg[63][7]  ( .D(n910), .E(n944), .CK(clk), .Q(\mem[63][7] ) );
  EDFFX1 \mem_reg[63][6]  ( .D(n905), .E(n944), .CK(clk), .Q(\mem[63][6] ) );
  EDFFX1 \mem_reg[63][5]  ( .D(n900), .E(n944), .CK(clk), .Q(\mem[63][5] ) );
  EDFFX1 \mem_reg[63][4]  ( .D(n895), .E(n944), .CK(clk), .Q(\mem[63][4] ) );
  EDFFX1 \mem_reg[63][3]  ( .D(n890), .E(n944), .CK(clk), .Q(\mem[63][3] ) );
  EDFFX1 \mem_reg[63][2]  ( .D(n885), .E(n944), .CK(clk), .Q(\mem[63][2] ) );
  EDFFX1 \mem_reg[63][1]  ( .D(n880), .E(n944), .CK(clk), .Q(\mem[63][1] ) );
  EDFFX1 \mem_reg[63][0]  ( .D(n875), .E(n944), .CK(clk), .Q(\mem[63][0] ) );
  EDFFX1 \mem_reg[67][7]  ( .D(n910), .E(n916), .CK(clk), .Q(\mem[67][7] ) );
  EDFFX1 \mem_reg[67][6]  ( .D(n905), .E(n916), .CK(clk), .Q(\mem[67][6] ) );
  EDFFX1 \mem_reg[67][5]  ( .D(n900), .E(n916), .CK(clk), .Q(\mem[67][5] ) );
  EDFFX1 \mem_reg[67][4]  ( .D(n895), .E(n916), .CK(clk), .Q(\mem[67][4] ) );
  EDFFX1 \mem_reg[67][3]  ( .D(n890), .E(n916), .CK(clk), .Q(\mem[67][3] ) );
  EDFFX1 \mem_reg[67][2]  ( .D(n885), .E(n916), .CK(clk), .Q(\mem[67][2] ) );
  EDFFX1 \mem_reg[67][1]  ( .D(n880), .E(n916), .CK(clk), .Q(\mem[67][1] ) );
  EDFFX1 \mem_reg[67][0]  ( .D(n875), .E(n916), .CK(clk), .Q(\mem[67][0] ) );
  EDFFX1 \mem_reg[71][7]  ( .D(n911), .E(n925), .CK(clk), .Q(\mem[71][7] ) );
  EDFFX1 \mem_reg[71][6]  ( .D(n906), .E(n925), .CK(clk), .Q(\mem[71][6] ) );
  EDFFX1 \mem_reg[71][5]  ( .D(n901), .E(n925), .CK(clk), .Q(\mem[71][5] ) );
  EDFFX1 \mem_reg[71][4]  ( .D(n896), .E(n925), .CK(clk), .Q(\mem[71][4] ) );
  EDFFX1 \mem_reg[71][3]  ( .D(n891), .E(n925), .CK(clk), .Q(\mem[71][3] ) );
  EDFFX1 \mem_reg[71][2]  ( .D(n886), .E(n925), .CK(clk), .Q(\mem[71][2] ) );
  EDFFX1 \mem_reg[71][1]  ( .D(n881), .E(n925), .CK(clk), .Q(\mem[71][1] ) );
  EDFFX1 \mem_reg[71][0]  ( .D(n876), .E(n925), .CK(clk), .Q(\mem[71][0] ) );
  EDFFX1 \mem_reg[75][7]  ( .D(n909), .E(n934), .CK(clk), .Q(\mem[75][7] ) );
  EDFFX1 \mem_reg[75][6]  ( .D(n904), .E(n934), .CK(clk), .Q(\mem[75][6] ) );
  EDFFX1 \mem_reg[75][5]  ( .D(n899), .E(n934), .CK(clk), .Q(\mem[75][5] ) );
  EDFFX1 \mem_reg[75][4]  ( .D(n894), .E(n934), .CK(clk), .Q(\mem[75][4] ) );
  EDFFX1 \mem_reg[75][3]  ( .D(n889), .E(n934), .CK(clk), .Q(\mem[75][3] ) );
  EDFFX1 \mem_reg[75][2]  ( .D(n884), .E(n934), .CK(clk), .Q(\mem[75][2] ) );
  EDFFX1 \mem_reg[75][1]  ( .D(n879), .E(n934), .CK(clk), .Q(\mem[75][1] ) );
  EDFFX1 \mem_reg[75][0]  ( .D(n874), .E(n934), .CK(clk), .Q(\mem[75][0] ) );
  EDFFX1 \mem_reg[79][7]  ( .D(n909), .E(n943), .CK(clk), .Q(\mem[79][7] ) );
  EDFFX1 \mem_reg[79][6]  ( .D(n904), .E(n943), .CK(clk), .Q(\mem[79][6] ) );
  EDFFX1 \mem_reg[79][5]  ( .D(n899), .E(n943), .CK(clk), .Q(\mem[79][5] ) );
  EDFFX1 \mem_reg[79][4]  ( .D(n894), .E(n943), .CK(clk), .Q(\mem[79][4] ) );
  EDFFX1 \mem_reg[79][3]  ( .D(n889), .E(n943), .CK(clk), .Q(\mem[79][3] ) );
  EDFFX1 \mem_reg[79][2]  ( .D(n884), .E(n943), .CK(clk), .Q(\mem[79][2] ) );
  EDFFX1 \mem_reg[79][1]  ( .D(n879), .E(n943), .CK(clk), .Q(\mem[79][1] ) );
  EDFFX1 \mem_reg[79][0]  ( .D(n874), .E(n943), .CK(clk), .Q(\mem[79][0] ) );
  EDFFX1 \mem_reg[83][7]  ( .D(n909), .E(n915), .CK(clk), .Q(\mem[83][7] ) );
  EDFFX1 \mem_reg[83][6]  ( .D(n904), .E(n915), .CK(clk), .Q(\mem[83][6] ) );
  EDFFX1 \mem_reg[83][5]  ( .D(n899), .E(n915), .CK(clk), .Q(\mem[83][5] ) );
  EDFFX1 \mem_reg[83][4]  ( .D(n894), .E(n915), .CK(clk), .Q(\mem[83][4] ) );
  EDFFX1 \mem_reg[83][3]  ( .D(n889), .E(n915), .CK(clk), .Q(\mem[83][3] ) );
  EDFFX1 \mem_reg[83][2]  ( .D(n884), .E(n915), .CK(clk), .Q(\mem[83][2] ) );
  EDFFX1 \mem_reg[83][1]  ( .D(n879), .E(n915), .CK(clk), .Q(\mem[83][1] ) );
  EDFFX1 \mem_reg[83][0]  ( .D(n874), .E(n915), .CK(clk), .Q(\mem[83][0] ) );
  EDFFX1 \mem_reg[87][7]  ( .D(n909), .E(n924), .CK(clk), .Q(\mem[87][7] ) );
  EDFFX1 \mem_reg[87][6]  ( .D(n904), .E(n924), .CK(clk), .Q(\mem[87][6] ) );
  EDFFX1 \mem_reg[87][5]  ( .D(n899), .E(n924), .CK(clk), .Q(\mem[87][5] ) );
  EDFFX1 \mem_reg[87][4]  ( .D(n894), .E(n924), .CK(clk), .Q(\mem[87][4] ) );
  EDFFX1 \mem_reg[87][3]  ( .D(n889), .E(n924), .CK(clk), .Q(\mem[87][3] ) );
  EDFFX1 \mem_reg[87][2]  ( .D(n884), .E(n924), .CK(clk), .Q(\mem[87][2] ) );
  EDFFX1 \mem_reg[87][1]  ( .D(n879), .E(n924), .CK(clk), .Q(\mem[87][1] ) );
  EDFFX1 \mem_reg[87][0]  ( .D(n874), .E(n924), .CK(clk), .Q(\mem[87][0] ) );
  EDFFX1 \mem_reg[91][7]  ( .D(n909), .E(n933), .CK(clk), .Q(\mem[91][7] ) );
  EDFFX1 \mem_reg[91][6]  ( .D(n904), .E(n933), .CK(clk), .Q(\mem[91][6] ) );
  EDFFX1 \mem_reg[91][5]  ( .D(n899), .E(n933), .CK(clk), .Q(\mem[91][5] ) );
  EDFFX1 \mem_reg[91][4]  ( .D(n894), .E(n933), .CK(clk), .Q(\mem[91][4] ) );
  EDFFX1 \mem_reg[91][3]  ( .D(n889), .E(n933), .CK(clk), .Q(\mem[91][3] ) );
  EDFFX1 \mem_reg[91][2]  ( .D(n884), .E(n933), .CK(clk), .Q(\mem[91][2] ) );
  EDFFX1 \mem_reg[91][1]  ( .D(n879), .E(n933), .CK(clk), .Q(\mem[91][1] ) );
  EDFFX1 \mem_reg[91][0]  ( .D(n874), .E(n933), .CK(clk), .Q(\mem[91][0] ) );
  EDFFX1 \mem_reg[95][7]  ( .D(n907), .E(n942), .CK(clk), .Q(\mem[95][7] ) );
  EDFFX1 \mem_reg[95][6]  ( .D(n902), .E(n942), .CK(clk), .Q(\mem[95][6] ) );
  EDFFX1 \mem_reg[95][5]  ( .D(n897), .E(n942), .CK(clk), .Q(\mem[95][5] ) );
  EDFFX1 \mem_reg[95][4]  ( .D(n892), .E(n942), .CK(clk), .Q(\mem[95][4] ) );
  EDFFX1 \mem_reg[95][3]  ( .D(n887), .E(n942), .CK(clk), .Q(\mem[95][3] ) );
  EDFFX1 \mem_reg[95][2]  ( .D(n882), .E(n942), .CK(clk), .Q(\mem[95][2] ) );
  EDFFX1 \mem_reg[95][1]  ( .D(n877), .E(n942), .CK(clk), .Q(\mem[95][1] ) );
  EDFFX1 \mem_reg[95][0]  ( .D(n872), .E(n942), .CK(clk), .Q(\mem[95][0] ) );
  EDFFX1 \mem_reg[99][7]  ( .D(n908), .E(n914), .CK(clk), .Q(\mem[99][7] ) );
  EDFFX1 \mem_reg[99][6]  ( .D(n903), .E(n914), .CK(clk), .Q(\mem[99][6] ) );
  EDFFX1 \mem_reg[99][5]  ( .D(n898), .E(n914), .CK(clk), .Q(\mem[99][5] ) );
  EDFFX1 \mem_reg[99][4]  ( .D(n893), .E(n914), .CK(clk), .Q(\mem[99][4] ) );
  EDFFX1 \mem_reg[99][3]  ( .D(n888), .E(n914), .CK(clk), .Q(\mem[99][3] ) );
  EDFFX1 \mem_reg[99][2]  ( .D(n883), .E(n914), .CK(clk), .Q(\mem[99][2] ) );
  EDFFX1 \mem_reg[99][1]  ( .D(n878), .E(n914), .CK(clk), .Q(\mem[99][1] ) );
  EDFFX1 \mem_reg[99][0]  ( .D(n873), .E(n914), .CK(clk), .Q(\mem[99][0] ) );
  EDFFX1 \mem_reg[103][7]  ( .D(n911), .E(n923), .CK(clk), .Q(\mem[103][7] )
         );
  EDFFX1 \mem_reg[103][6]  ( .D(n906), .E(n923), .CK(clk), .Q(\mem[103][6] )
         );
  EDFFX1 \mem_reg[103][5]  ( .D(n901), .E(n923), .CK(clk), .Q(\mem[103][5] )
         );
  EDFFX1 \mem_reg[103][4]  ( .D(n896), .E(n923), .CK(clk), .Q(\mem[103][4] )
         );
  EDFFX1 \mem_reg[103][3]  ( .D(n891), .E(n923), .CK(clk), .Q(\mem[103][3] )
         );
  EDFFX1 \mem_reg[103][2]  ( .D(n886), .E(n923), .CK(clk), .Q(\mem[103][2] )
         );
  EDFFX1 \mem_reg[103][1]  ( .D(n881), .E(n923), .CK(clk), .Q(\mem[103][1] )
         );
  EDFFX1 \mem_reg[103][0]  ( .D(n876), .E(n923), .CK(clk), .Q(\mem[103][0] )
         );
  EDFFX1 \mem_reg[107][7]  ( .D(n908), .E(n932), .CK(clk), .Q(\mem[107][7] )
         );
  EDFFX1 \mem_reg[107][6]  ( .D(n903), .E(n932), .CK(clk), .Q(\mem[107][6] )
         );
  EDFFX1 \mem_reg[107][5]  ( .D(n898), .E(n932), .CK(clk), .Q(\mem[107][5] )
         );
  EDFFX1 \mem_reg[107][4]  ( .D(n893), .E(n932), .CK(clk), .Q(\mem[107][4] )
         );
  EDFFX1 \mem_reg[107][3]  ( .D(n888), .E(n932), .CK(clk), .Q(\mem[107][3] )
         );
  EDFFX1 \mem_reg[107][2]  ( .D(n883), .E(n932), .CK(clk), .Q(\mem[107][2] )
         );
  EDFFX1 \mem_reg[107][1]  ( .D(n878), .E(n932), .CK(clk), .Q(\mem[107][1] )
         );
  EDFFX1 \mem_reg[107][0]  ( .D(n873), .E(n932), .CK(clk), .Q(\mem[107][0] )
         );
  EDFFX1 \mem_reg[111][7]  ( .D(n908), .E(n941), .CK(clk), .Q(\mem[111][7] )
         );
  EDFFX1 \mem_reg[111][6]  ( .D(n903), .E(n941), .CK(clk), .Q(\mem[111][6] )
         );
  EDFFX1 \mem_reg[111][5]  ( .D(n898), .E(n941), .CK(clk), .Q(\mem[111][5] )
         );
  EDFFX1 \mem_reg[111][4]  ( .D(n893), .E(n941), .CK(clk), .Q(\mem[111][4] )
         );
  EDFFX1 \mem_reg[111][3]  ( .D(n888), .E(n941), .CK(clk), .Q(\mem[111][3] )
         );
  EDFFX1 \mem_reg[111][2]  ( .D(n883), .E(n941), .CK(clk), .Q(\mem[111][2] )
         );
  EDFFX1 \mem_reg[111][1]  ( .D(n878), .E(n941), .CK(clk), .Q(\mem[111][1] )
         );
  EDFFX1 \mem_reg[111][0]  ( .D(n873), .E(n941), .CK(clk), .Q(\mem[111][0] )
         );
  EDFFX1 \mem_reg[115][7]  ( .D(n908), .E(n913), .CK(clk), .Q(\mem[115][7] )
         );
  EDFFX1 \mem_reg[115][6]  ( .D(n903), .E(n913), .CK(clk), .Q(\mem[115][6] )
         );
  EDFFX1 \mem_reg[115][5]  ( .D(n898), .E(n913), .CK(clk), .Q(\mem[115][5] )
         );
  EDFFX1 \mem_reg[115][4]  ( .D(n893), .E(n913), .CK(clk), .Q(\mem[115][4] )
         );
  EDFFX1 \mem_reg[115][3]  ( .D(n888), .E(n913), .CK(clk), .Q(\mem[115][3] )
         );
  EDFFX1 \mem_reg[115][2]  ( .D(n883), .E(n913), .CK(clk), .Q(\mem[115][2] )
         );
  EDFFX1 \mem_reg[115][1]  ( .D(n878), .E(n913), .CK(clk), .Q(\mem[115][1] )
         );
  EDFFX1 \mem_reg[115][0]  ( .D(n873), .E(n913), .CK(clk), .Q(\mem[115][0] )
         );
  EDFFX1 \mem_reg[119][7]  ( .D(n907), .E(n922), .CK(clk), .Q(\mem[119][7] )
         );
  EDFFX1 \mem_reg[119][6]  ( .D(n902), .E(n922), .CK(clk), .Q(\mem[119][6] )
         );
  EDFFX1 \mem_reg[119][5]  ( .D(n897), .E(n922), .CK(clk), .Q(\mem[119][5] )
         );
  EDFFX1 \mem_reg[119][4]  ( .D(n892), .E(n922), .CK(clk), .Q(\mem[119][4] )
         );
  EDFFX1 \mem_reg[119][3]  ( .D(n887), .E(n922), .CK(clk), .Q(\mem[119][3] )
         );
  EDFFX1 \mem_reg[119][2]  ( .D(n882), .E(n922), .CK(clk), .Q(\mem[119][2] )
         );
  EDFFX1 \mem_reg[119][1]  ( .D(n877), .E(n922), .CK(clk), .Q(\mem[119][1] )
         );
  EDFFX1 \mem_reg[119][0]  ( .D(n872), .E(n922), .CK(clk), .Q(\mem[119][0] )
         );
  EDFFX1 \mem_reg[123][7]  ( .D(n907), .E(n931), .CK(clk), .Q(\mem[123][7] )
         );
  EDFFX1 \mem_reg[123][6]  ( .D(n902), .E(n931), .CK(clk), .Q(\mem[123][6] )
         );
  EDFFX1 \mem_reg[123][5]  ( .D(n897), .E(n931), .CK(clk), .Q(\mem[123][5] )
         );
  EDFFX1 \mem_reg[123][4]  ( .D(n892), .E(n931), .CK(clk), .Q(\mem[123][4] )
         );
  EDFFX1 \mem_reg[123][3]  ( .D(n887), .E(n931), .CK(clk), .Q(\mem[123][3] )
         );
  EDFFX1 \mem_reg[123][2]  ( .D(n882), .E(n931), .CK(clk), .Q(\mem[123][2] )
         );
  EDFFX1 \mem_reg[123][1]  ( .D(n877), .E(n931), .CK(clk), .Q(\mem[123][1] )
         );
  EDFFX1 \mem_reg[123][0]  ( .D(n872), .E(n931), .CK(clk), .Q(\mem[123][0] )
         );
  EDFFX1 \mem_reg[127][7]  ( .D(n907), .E(n940), .CK(clk), .Q(\mem[127][7] )
         );
  EDFFX1 \mem_reg[127][6]  ( .D(n902), .E(n940), .CK(clk), .Q(\mem[127][6] )
         );
  EDFFX1 \mem_reg[127][5]  ( .D(n897), .E(n940), .CK(clk), .Q(\mem[127][5] )
         );
  EDFFX1 \mem_reg[127][4]  ( .D(n892), .E(n940), .CK(clk), .Q(\mem[127][4] )
         );
  EDFFX1 \mem_reg[127][3]  ( .D(n887), .E(n940), .CK(clk), .Q(\mem[127][3] )
         );
  EDFFX1 \mem_reg[127][2]  ( .D(n882), .E(n940), .CK(clk), .Q(\mem[127][2] )
         );
  EDFFX1 \mem_reg[127][1]  ( .D(n877), .E(n940), .CK(clk), .Q(\mem[127][1] )
         );
  EDFFX1 \mem_reg[127][0]  ( .D(n872), .E(n940), .CK(clk), .Q(\mem[127][0] )
         );
  EDFFX1 \mem_reg[0][7]  ( .D(n907), .E(n993), .CK(clk), .Q(\mem[0][7] ) );
  EDFFX1 \mem_reg[0][6]  ( .D(n902), .E(n993), .CK(clk), .Q(\mem[0][6] ) );
  EDFFX1 \mem_reg[0][5]  ( .D(n897), .E(n993), .CK(clk), .Q(\mem[0][5] ) );
  EDFFX1 \mem_reg[0][4]  ( .D(n892), .E(n993), .CK(clk), .Q(\mem[0][4] ) );
  EDFFX1 \mem_reg[0][3]  ( .D(n887), .E(n993), .CK(clk), .Q(\mem[0][3] ) );
  EDFFX1 \mem_reg[0][2]  ( .D(n882), .E(n993), .CK(clk), .Q(\mem[0][2] ) );
  EDFFX1 \mem_reg[0][1]  ( .D(n877), .E(n993), .CK(clk), .Q(\mem[0][1] ) );
  EDFFX1 \mem_reg[0][0]  ( .D(n872), .E(n993), .CK(clk), .Q(\mem[0][0] ) );
  EDFFX1 \mem_reg[4][7]  ( .D(n908), .E(n1002), .CK(clk), .Q(\mem[4][7] ) );
  EDFFX1 \mem_reg[4][6]  ( .D(n903), .E(n1002), .CK(clk), .Q(\mem[4][6] ) );
  EDFFX1 \mem_reg[4][5]  ( .D(n898), .E(n1002), .CK(clk), .Q(\mem[4][5] ) );
  EDFFX1 \mem_reg[4][4]  ( .D(n893), .E(n1002), .CK(clk), .Q(\mem[4][4] ) );
  EDFFX1 \mem_reg[4][3]  ( .D(n888), .E(n1002), .CK(clk), .Q(\mem[4][3] ) );
  EDFFX1 \mem_reg[4][2]  ( .D(n883), .E(n1002), .CK(clk), .Q(\mem[4][2] ) );
  EDFFX1 \mem_reg[4][1]  ( .D(n878), .E(n1002), .CK(clk), .Q(\mem[4][1] ) );
  EDFFX1 \mem_reg[4][0]  ( .D(n873), .E(n1002), .CK(clk), .Q(\mem[4][0] ) );
  EDFFX1 \mem_reg[8][7]  ( .D(n911), .E(n1011), .CK(clk), .Q(\mem[8][7] ) );
  EDFFX1 \mem_reg[8][6]  ( .D(n906), .E(n1011), .CK(clk), .Q(\mem[8][6] ) );
  EDFFX1 \mem_reg[8][5]  ( .D(n901), .E(n1011), .CK(clk), .Q(\mem[8][5] ) );
  EDFFX1 \mem_reg[8][4]  ( .D(n896), .E(n1011), .CK(clk), .Q(\mem[8][4] ) );
  EDFFX1 \mem_reg[8][3]  ( .D(n891), .E(n1011), .CK(clk), .Q(\mem[8][3] ) );
  EDFFX1 \mem_reg[8][2]  ( .D(n886), .E(n1011), .CK(clk), .Q(\mem[8][2] ) );
  EDFFX1 \mem_reg[8][1]  ( .D(n881), .E(n1011), .CK(clk), .Q(\mem[8][1] ) );
  EDFFX1 \mem_reg[8][0]  ( .D(n876), .E(n1011), .CK(clk), .Q(\mem[8][0] ) );
  EDFFX1 \mem_reg[12][7]  ( .D(n910), .E(n1020), .CK(clk), .Q(\mem[12][7] ) );
  EDFFX1 \mem_reg[12][6]  ( .D(n905), .E(n1020), .CK(clk), .Q(\mem[12][6] ) );
  EDFFX1 \mem_reg[12][5]  ( .D(n900), .E(n1020), .CK(clk), .Q(\mem[12][5] ) );
  EDFFX1 \mem_reg[12][4]  ( .D(n895), .E(n1020), .CK(clk), .Q(\mem[12][4] ) );
  EDFFX1 \mem_reg[12][3]  ( .D(n890), .E(n1020), .CK(clk), .Q(\mem[12][3] ) );
  EDFFX1 \mem_reg[12][2]  ( .D(n885), .E(n1020), .CK(clk), .Q(\mem[12][2] ) );
  EDFFX1 \mem_reg[12][1]  ( .D(n880), .E(n1020), .CK(clk), .Q(\mem[12][1] ) );
  EDFFX1 \mem_reg[12][0]  ( .D(n875), .E(n1020), .CK(clk), .Q(\mem[12][0] ) );
  EDFFX1 \mem_reg[16][7]  ( .D(n910), .E(n992), .CK(clk), .Q(\mem[16][7] ) );
  EDFFX1 \mem_reg[16][6]  ( .D(n905), .E(n992), .CK(clk), .Q(\mem[16][6] ) );
  EDFFX1 \mem_reg[16][5]  ( .D(n900), .E(n992), .CK(clk), .Q(\mem[16][5] ) );
  EDFFX1 \mem_reg[16][4]  ( .D(n895), .E(n992), .CK(clk), .Q(\mem[16][4] ) );
  EDFFX1 \mem_reg[16][3]  ( .D(n890), .E(n992), .CK(clk), .Q(\mem[16][3] ) );
  EDFFX1 \mem_reg[16][2]  ( .D(n885), .E(n992), .CK(clk), .Q(\mem[16][2] ) );
  EDFFX1 \mem_reg[16][1]  ( .D(n880), .E(n992), .CK(clk), .Q(\mem[16][1] ) );
  EDFFX1 \mem_reg[16][0]  ( .D(n875), .E(n992), .CK(clk), .Q(\mem[16][0] ) );
  EDFFX1 \mem_reg[20][7]  ( .D(data_in[7]), .E(n1001), .CK(clk), .Q(
        \mem[20][7] ) );
  EDFFX1 \mem_reg[20][6]  ( .D(data_in[6]), .E(n1001), .CK(clk), .Q(
        \mem[20][6] ) );
  EDFFX1 \mem_reg[20][5]  ( .D(data_in[5]), .E(n1001), .CK(clk), .Q(
        \mem[20][5] ) );
  EDFFX1 \mem_reg[20][4]  ( .D(data_in[4]), .E(n1001), .CK(clk), .Q(
        \mem[20][4] ) );
  EDFFX1 \mem_reg[20][3]  ( .D(data_in[3]), .E(n1001), .CK(clk), .Q(
        \mem[20][3] ) );
  EDFFX1 \mem_reg[20][2]  ( .D(data_in[2]), .E(n1001), .CK(clk), .Q(
        \mem[20][2] ) );
  EDFFX1 \mem_reg[20][1]  ( .D(data_in[1]), .E(n1001), .CK(clk), .Q(
        \mem[20][1] ) );
  EDFFX1 \mem_reg[20][0]  ( .D(data_in[0]), .E(n1001), .CK(clk), .Q(
        \mem[20][0] ) );
  EDFFX1 \mem_reg[24][7]  ( .D(data_in[7]), .E(n1010), .CK(clk), .Q(
        \mem[24][7] ) );
  EDFFX1 \mem_reg[24][6]  ( .D(data_in[6]), .E(n1010), .CK(clk), .Q(
        \mem[24][6] ) );
  EDFFX1 \mem_reg[24][5]  ( .D(data_in[5]), .E(n1010), .CK(clk), .Q(
        \mem[24][5] ) );
  EDFFX1 \mem_reg[24][4]  ( .D(data_in[4]), .E(n1010), .CK(clk), .Q(
        \mem[24][4] ) );
  EDFFX1 \mem_reg[24][3]  ( .D(data_in[3]), .E(n1010), .CK(clk), .Q(
        \mem[24][3] ) );
  EDFFX1 \mem_reg[24][2]  ( .D(data_in[2]), .E(n1010), .CK(clk), .Q(
        \mem[24][2] ) );
  EDFFX1 \mem_reg[24][1]  ( .D(data_in[1]), .E(n1010), .CK(clk), .Q(
        \mem[24][1] ) );
  EDFFX1 \mem_reg[24][0]  ( .D(data_in[0]), .E(n1010), .CK(clk), .Q(
        \mem[24][0] ) );
  EDFFX1 \mem_reg[28][7]  ( .D(data_in[7]), .E(n1019), .CK(clk), .Q(
        \mem[28][7] ) );
  EDFFX1 \mem_reg[28][6]  ( .D(data_in[6]), .E(n1019), .CK(clk), .Q(
        \mem[28][6] ) );
  EDFFX1 \mem_reg[28][5]  ( .D(data_in[5]), .E(n1019), .CK(clk), .Q(
        \mem[28][5] ) );
  EDFFX1 \mem_reg[28][4]  ( .D(data_in[4]), .E(n1019), .CK(clk), .Q(
        \mem[28][4] ) );
  EDFFX1 \mem_reg[28][3]  ( .D(data_in[3]), .E(n1019), .CK(clk), .Q(
        \mem[28][3] ) );
  EDFFX1 \mem_reg[28][2]  ( .D(data_in[2]), .E(n1019), .CK(clk), .Q(
        \mem[28][2] ) );
  EDFFX1 \mem_reg[28][1]  ( .D(data_in[1]), .E(n1019), .CK(clk), .Q(
        \mem[28][1] ) );
  EDFFX1 \mem_reg[28][0]  ( .D(data_in[0]), .E(n1019), .CK(clk), .Q(
        \mem[28][0] ) );
  EDFFX1 \mem_reg[32][7]  ( .D(n911), .E(n991), .CK(clk), .Q(\mem[32][7] ) );
  EDFFX1 \mem_reg[32][6]  ( .D(n906), .E(n991), .CK(clk), .Q(\mem[32][6] ) );
  EDFFX1 \mem_reg[32][5]  ( .D(n901), .E(n991), .CK(clk), .Q(\mem[32][5] ) );
  EDFFX1 \mem_reg[32][4]  ( .D(n896), .E(n991), .CK(clk), .Q(\mem[32][4] ) );
  EDFFX1 \mem_reg[32][3]  ( .D(n891), .E(n991), .CK(clk), .Q(\mem[32][3] ) );
  EDFFX1 \mem_reg[32][2]  ( .D(n886), .E(n991), .CK(clk), .Q(\mem[32][2] ) );
  EDFFX1 \mem_reg[32][1]  ( .D(n881), .E(n991), .CK(clk), .Q(\mem[32][1] ) );
  EDFFX1 \mem_reg[32][0]  ( .D(n876), .E(n991), .CK(clk), .Q(\mem[32][0] ) );
  EDFFX1 \mem_reg[36][7]  ( .D(n911), .E(n1000), .CK(clk), .Q(\mem[36][7] ) );
  EDFFX1 \mem_reg[36][6]  ( .D(n906), .E(n1000), .CK(clk), .Q(\mem[36][6] ) );
  EDFFX1 \mem_reg[36][5]  ( .D(n901), .E(n1000), .CK(clk), .Q(\mem[36][5] ) );
  EDFFX1 \mem_reg[36][4]  ( .D(n896), .E(n1000), .CK(clk), .Q(\mem[36][4] ) );
  EDFFX1 \mem_reg[36][3]  ( .D(n891), .E(n1000), .CK(clk), .Q(\mem[36][3] ) );
  EDFFX1 \mem_reg[36][2]  ( .D(n886), .E(n1000), .CK(clk), .Q(\mem[36][2] ) );
  EDFFX1 \mem_reg[36][1]  ( .D(n881), .E(n1000), .CK(clk), .Q(\mem[36][1] ) );
  EDFFX1 \mem_reg[36][0]  ( .D(n876), .E(n1000), .CK(clk), .Q(\mem[36][0] ) );
  EDFFX1 \mem_reg[40][7]  ( .D(n911), .E(n1009), .CK(clk), .Q(\mem[40][7] ) );
  EDFFX1 \mem_reg[40][6]  ( .D(n906), .E(n1009), .CK(clk), .Q(\mem[40][6] ) );
  EDFFX1 \mem_reg[40][5]  ( .D(n901), .E(n1009), .CK(clk), .Q(\mem[40][5] ) );
  EDFFX1 \mem_reg[40][4]  ( .D(n896), .E(n1009), .CK(clk), .Q(\mem[40][4] ) );
  EDFFX1 \mem_reg[40][3]  ( .D(n891), .E(n1009), .CK(clk), .Q(\mem[40][3] ) );
  EDFFX1 \mem_reg[40][2]  ( .D(n886), .E(n1009), .CK(clk), .Q(\mem[40][2] ) );
  EDFFX1 \mem_reg[40][1]  ( .D(n881), .E(n1009), .CK(clk), .Q(\mem[40][1] ) );
  EDFFX1 \mem_reg[40][0]  ( .D(n876), .E(n1009), .CK(clk), .Q(\mem[40][0] ) );
  EDFFX1 \mem_reg[44][7]  ( .D(n910), .E(n1018), .CK(clk), .Q(\mem[44][7] ) );
  EDFFX1 \mem_reg[44][6]  ( .D(n905), .E(n1018), .CK(clk), .Q(\mem[44][6] ) );
  EDFFX1 \mem_reg[44][5]  ( .D(n900), .E(n1018), .CK(clk), .Q(\mem[44][5] ) );
  EDFFX1 \mem_reg[44][4]  ( .D(n895), .E(n1018), .CK(clk), .Q(\mem[44][4] ) );
  EDFFX1 \mem_reg[44][3]  ( .D(n890), .E(n1018), .CK(clk), .Q(\mem[44][3] ) );
  EDFFX1 \mem_reg[44][2]  ( .D(n885), .E(n1018), .CK(clk), .Q(\mem[44][2] ) );
  EDFFX1 \mem_reg[44][1]  ( .D(n880), .E(n1018), .CK(clk), .Q(\mem[44][1] ) );
  EDFFX1 \mem_reg[44][0]  ( .D(n875), .E(n1018), .CK(clk), .Q(\mem[44][0] ) );
  EDFFX1 \mem_reg[48][7]  ( .D(n907), .E(n990), .CK(clk), .Q(\mem[48][7] ) );
  EDFFX1 \mem_reg[48][6]  ( .D(n902), .E(n990), .CK(clk), .Q(\mem[48][6] ) );
  EDFFX1 \mem_reg[48][5]  ( .D(n897), .E(n990), .CK(clk), .Q(\mem[48][5] ) );
  EDFFX1 \mem_reg[48][4]  ( .D(n892), .E(n990), .CK(clk), .Q(\mem[48][4] ) );
  EDFFX1 \mem_reg[48][3]  ( .D(n887), .E(n990), .CK(clk), .Q(\mem[48][3] ) );
  EDFFX1 \mem_reg[48][2]  ( .D(n882), .E(n990), .CK(clk), .Q(\mem[48][2] ) );
  EDFFX1 \mem_reg[48][1]  ( .D(n877), .E(n990), .CK(clk), .Q(\mem[48][1] ) );
  EDFFX1 \mem_reg[48][0]  ( .D(n872), .E(n990), .CK(clk), .Q(\mem[48][0] ) );
  EDFFX1 \mem_reg[52][7]  ( .D(n908), .E(n999), .CK(clk), .Q(\mem[52][7] ) );
  EDFFX1 \mem_reg[52][6]  ( .D(n903), .E(n999), .CK(clk), .Q(\mem[52][6] ) );
  EDFFX1 \mem_reg[52][5]  ( .D(n898), .E(n999), .CK(clk), .Q(\mem[52][5] ) );
  EDFFX1 \mem_reg[52][4]  ( .D(n893), .E(n999), .CK(clk), .Q(\mem[52][4] ) );
  EDFFX1 \mem_reg[52][3]  ( .D(n888), .E(n999), .CK(clk), .Q(\mem[52][3] ) );
  EDFFX1 \mem_reg[52][2]  ( .D(n883), .E(n999), .CK(clk), .Q(\mem[52][2] ) );
  EDFFX1 \mem_reg[52][1]  ( .D(n878), .E(n999), .CK(clk), .Q(\mem[52][1] ) );
  EDFFX1 \mem_reg[52][0]  ( .D(n873), .E(n999), .CK(clk), .Q(\mem[52][0] ) );
  EDFFX1 \mem_reg[56][7]  ( .D(n910), .E(n1008), .CK(clk), .Q(\mem[56][7] ) );
  EDFFX1 \mem_reg[56][6]  ( .D(n905), .E(n1008), .CK(clk), .Q(\mem[56][6] ) );
  EDFFX1 \mem_reg[56][5]  ( .D(n900), .E(n1008), .CK(clk), .Q(\mem[56][5] ) );
  EDFFX1 \mem_reg[56][4]  ( .D(n895), .E(n1008), .CK(clk), .Q(\mem[56][4] ) );
  EDFFX1 \mem_reg[56][3]  ( .D(n890), .E(n1008), .CK(clk), .Q(\mem[56][3] ) );
  EDFFX1 \mem_reg[56][2]  ( .D(n885), .E(n1008), .CK(clk), .Q(\mem[56][2] ) );
  EDFFX1 \mem_reg[56][1]  ( .D(n880), .E(n1008), .CK(clk), .Q(\mem[56][1] ) );
  EDFFX1 \mem_reg[56][0]  ( .D(n875), .E(n1008), .CK(clk), .Q(\mem[56][0] ) );
  EDFFX1 \mem_reg[60][7]  ( .D(n910), .E(n1017), .CK(clk), .Q(\mem[60][7] ) );
  EDFFX1 \mem_reg[60][6]  ( .D(n905), .E(n1017), .CK(clk), .Q(\mem[60][6] ) );
  EDFFX1 \mem_reg[60][5]  ( .D(n900), .E(n1017), .CK(clk), .Q(\mem[60][5] ) );
  EDFFX1 \mem_reg[60][4]  ( .D(n895), .E(n1017), .CK(clk), .Q(\mem[60][4] ) );
  EDFFX1 \mem_reg[60][3]  ( .D(n890), .E(n1017), .CK(clk), .Q(\mem[60][3] ) );
  EDFFX1 \mem_reg[60][2]  ( .D(n885), .E(n1017), .CK(clk), .Q(\mem[60][2] ) );
  EDFFX1 \mem_reg[60][1]  ( .D(n880), .E(n1017), .CK(clk), .Q(\mem[60][1] ) );
  EDFFX1 \mem_reg[60][0]  ( .D(n875), .E(n1017), .CK(clk), .Q(\mem[60][0] ) );
  EDFFX1 \mem_reg[64][7]  ( .D(n910), .E(n989), .CK(clk), .Q(\mem[64][7] ) );
  EDFFX1 \mem_reg[64][6]  ( .D(n905), .E(n989), .CK(clk), .Q(\mem[64][6] ) );
  EDFFX1 \mem_reg[64][5]  ( .D(n900), .E(n989), .CK(clk), .Q(\mem[64][5] ) );
  EDFFX1 \mem_reg[64][4]  ( .D(n895), .E(n989), .CK(clk), .Q(\mem[64][4] ) );
  EDFFX1 \mem_reg[64][3]  ( .D(n890), .E(n989), .CK(clk), .Q(\mem[64][3] ) );
  EDFFX1 \mem_reg[64][2]  ( .D(n885), .E(n989), .CK(clk), .Q(\mem[64][2] ) );
  EDFFX1 \mem_reg[64][1]  ( .D(n880), .E(n989), .CK(clk), .Q(\mem[64][1] ) );
  EDFFX1 \mem_reg[64][0]  ( .D(n875), .E(n989), .CK(clk), .Q(\mem[64][0] ) );
  EDFFX1 \mem_reg[68][7]  ( .D(n909), .E(n998), .CK(clk), .Q(\mem[68][7] ) );
  EDFFX1 \mem_reg[68][6]  ( .D(n904), .E(n998), .CK(clk), .Q(\mem[68][6] ) );
  EDFFX1 \mem_reg[68][5]  ( .D(n899), .E(n998), .CK(clk), .Q(\mem[68][5] ) );
  EDFFX1 \mem_reg[68][4]  ( .D(n894), .E(n998), .CK(clk), .Q(\mem[68][4] ) );
  EDFFX1 \mem_reg[68][3]  ( .D(n889), .E(n998), .CK(clk), .Q(\mem[68][3] ) );
  EDFFX1 \mem_reg[68][2]  ( .D(n884), .E(n998), .CK(clk), .Q(\mem[68][2] ) );
  EDFFX1 \mem_reg[68][1]  ( .D(n879), .E(n998), .CK(clk), .Q(\mem[68][1] ) );
  EDFFX1 \mem_reg[68][0]  ( .D(n874), .E(n998), .CK(clk), .Q(\mem[68][0] ) );
  EDFFX1 \mem_reg[72][7]  ( .D(n909), .E(n1007), .CK(clk), .Q(\mem[72][7] ) );
  EDFFX1 \mem_reg[72][6]  ( .D(n904), .E(n1007), .CK(clk), .Q(\mem[72][6] ) );
  EDFFX1 \mem_reg[72][5]  ( .D(n899), .E(n1007), .CK(clk), .Q(\mem[72][5] ) );
  EDFFX1 \mem_reg[72][4]  ( .D(n894), .E(n1007), .CK(clk), .Q(\mem[72][4] ) );
  EDFFX1 \mem_reg[72][3]  ( .D(n889), .E(n1007), .CK(clk), .Q(\mem[72][3] ) );
  EDFFX1 \mem_reg[72][2]  ( .D(n884), .E(n1007), .CK(clk), .Q(\mem[72][2] ) );
  EDFFX1 \mem_reg[72][1]  ( .D(n879), .E(n1007), .CK(clk), .Q(\mem[72][1] ) );
  EDFFX1 \mem_reg[72][0]  ( .D(n874), .E(n1007), .CK(clk), .Q(\mem[72][0] ) );
  EDFFX1 \mem_reg[76][7]  ( .D(n909), .E(n1016), .CK(clk), .Q(\mem[76][7] ) );
  EDFFX1 \mem_reg[76][6]  ( .D(n904), .E(n1016), .CK(clk), .Q(\mem[76][6] ) );
  EDFFX1 \mem_reg[76][5]  ( .D(n899), .E(n1016), .CK(clk), .Q(\mem[76][5] ) );
  EDFFX1 \mem_reg[76][4]  ( .D(n894), .E(n1016), .CK(clk), .Q(\mem[76][4] ) );
  EDFFX1 \mem_reg[76][3]  ( .D(n889), .E(n1016), .CK(clk), .Q(\mem[76][3] ) );
  EDFFX1 \mem_reg[76][2]  ( .D(n884), .E(n1016), .CK(clk), .Q(\mem[76][2] ) );
  EDFFX1 \mem_reg[76][1]  ( .D(n879), .E(n1016), .CK(clk), .Q(\mem[76][1] ) );
  EDFFX1 \mem_reg[76][0]  ( .D(n874), .E(n1016), .CK(clk), .Q(\mem[76][0] ) );
  EDFFX1 \mem_reg[80][7]  ( .D(n909), .E(n988), .CK(clk), .Q(\mem[80][7] ) );
  EDFFX1 \mem_reg[80][6]  ( .D(n904), .E(n988), .CK(clk), .Q(\mem[80][6] ) );
  EDFFX1 \mem_reg[80][5]  ( .D(n899), .E(n988), .CK(clk), .Q(\mem[80][5] ) );
  EDFFX1 \mem_reg[80][4]  ( .D(n894), .E(n988), .CK(clk), .Q(\mem[80][4] ) );
  EDFFX1 \mem_reg[80][3]  ( .D(n889), .E(n988), .CK(clk), .Q(\mem[80][3] ) );
  EDFFX1 \mem_reg[80][2]  ( .D(n884), .E(n988), .CK(clk), .Q(\mem[80][2] ) );
  EDFFX1 \mem_reg[80][1]  ( .D(n879), .E(n988), .CK(clk), .Q(\mem[80][1] ) );
  EDFFX1 \mem_reg[80][0]  ( .D(n874), .E(n988), .CK(clk), .Q(\mem[80][0] ) );
  EDFFX1 \mem_reg[84][7]  ( .D(n909), .E(n997), .CK(clk), .Q(\mem[84][7] ) );
  EDFFX1 \mem_reg[84][6]  ( .D(n904), .E(n997), .CK(clk), .Q(\mem[84][6] ) );
  EDFFX1 \mem_reg[84][5]  ( .D(n899), .E(n997), .CK(clk), .Q(\mem[84][5] ) );
  EDFFX1 \mem_reg[84][4]  ( .D(n894), .E(n997), .CK(clk), .Q(\mem[84][4] ) );
  EDFFX1 \mem_reg[84][3]  ( .D(n889), .E(n997), .CK(clk), .Q(\mem[84][3] ) );
  EDFFX1 \mem_reg[84][2]  ( .D(n884), .E(n997), .CK(clk), .Q(\mem[84][2] ) );
  EDFFX1 \mem_reg[84][1]  ( .D(n879), .E(n997), .CK(clk), .Q(\mem[84][1] ) );
  EDFFX1 \mem_reg[84][0]  ( .D(n874), .E(n997), .CK(clk), .Q(\mem[84][0] ) );
  EDFFX1 \mem_reg[88][7]  ( .D(n909), .E(n1006), .CK(clk), .Q(\mem[88][7] ) );
  EDFFX1 \mem_reg[88][6]  ( .D(n904), .E(n1006), .CK(clk), .Q(\mem[88][6] ) );
  EDFFX1 \mem_reg[88][5]  ( .D(n899), .E(n1006), .CK(clk), .Q(\mem[88][5] ) );
  EDFFX1 \mem_reg[88][4]  ( .D(n894), .E(n1006), .CK(clk), .Q(\mem[88][4] ) );
  EDFFX1 \mem_reg[88][3]  ( .D(n889), .E(n1006), .CK(clk), .Q(\mem[88][3] ) );
  EDFFX1 \mem_reg[88][2]  ( .D(n884), .E(n1006), .CK(clk), .Q(\mem[88][2] ) );
  EDFFX1 \mem_reg[88][1]  ( .D(n879), .E(n1006), .CK(clk), .Q(\mem[88][1] ) );
  EDFFX1 \mem_reg[88][0]  ( .D(n874), .E(n1006), .CK(clk), .Q(\mem[88][0] ) );
  EDFFX1 \mem_reg[92][7]  ( .D(n911), .E(n1015), .CK(clk), .Q(\mem[92][7] ) );
  EDFFX1 \mem_reg[92][6]  ( .D(n906), .E(n1015), .CK(clk), .Q(\mem[92][6] ) );
  EDFFX1 \mem_reg[92][5]  ( .D(n901), .E(n1015), .CK(clk), .Q(\mem[92][5] ) );
  EDFFX1 \mem_reg[92][4]  ( .D(n896), .E(n1015), .CK(clk), .Q(\mem[92][4] ) );
  EDFFX1 \mem_reg[92][3]  ( .D(n891), .E(n1015), .CK(clk), .Q(\mem[92][3] ) );
  EDFFX1 \mem_reg[92][2]  ( .D(n886), .E(n1015), .CK(clk), .Q(\mem[92][2] ) );
  EDFFX1 \mem_reg[92][1]  ( .D(n881), .E(n1015), .CK(clk), .Q(\mem[92][1] ) );
  EDFFX1 \mem_reg[92][0]  ( .D(n876), .E(n1015), .CK(clk), .Q(\mem[92][0] ) );
  EDFFX1 \mem_reg[96][7]  ( .D(n910), .E(n987), .CK(clk), .Q(\mem[96][7] ) );
  EDFFX1 \mem_reg[96][6]  ( .D(n905), .E(n987), .CK(clk), .Q(\mem[96][6] ) );
  EDFFX1 \mem_reg[96][5]  ( .D(n900), .E(n987), .CK(clk), .Q(\mem[96][5] ) );
  EDFFX1 \mem_reg[96][4]  ( .D(n895), .E(n987), .CK(clk), .Q(\mem[96][4] ) );
  EDFFX1 \mem_reg[96][3]  ( .D(n890), .E(n987), .CK(clk), .Q(\mem[96][3] ) );
  EDFFX1 \mem_reg[96][2]  ( .D(n885), .E(n987), .CK(clk), .Q(\mem[96][2] ) );
  EDFFX1 \mem_reg[96][1]  ( .D(n880), .E(n987), .CK(clk), .Q(\mem[96][1] ) );
  EDFFX1 \mem_reg[96][0]  ( .D(n875), .E(n987), .CK(clk), .Q(\mem[96][0] ) );
  EDFFX1 \mem_reg[100][7]  ( .D(n907), .E(n996), .CK(clk), .Q(\mem[100][7] )
         );
  EDFFX1 \mem_reg[100][6]  ( .D(n902), .E(n996), .CK(clk), .Q(\mem[100][6] )
         );
  EDFFX1 \mem_reg[100][5]  ( .D(n897), .E(n996), .CK(clk), .Q(\mem[100][5] )
         );
  EDFFX1 \mem_reg[100][4]  ( .D(n892), .E(n996), .CK(clk), .Q(\mem[100][4] )
         );
  EDFFX1 \mem_reg[100][3]  ( .D(n887), .E(n996), .CK(clk), .Q(\mem[100][3] )
         );
  EDFFX1 \mem_reg[100][2]  ( .D(n882), .E(n996), .CK(clk), .Q(\mem[100][2] )
         );
  EDFFX1 \mem_reg[100][1]  ( .D(n877), .E(n996), .CK(clk), .Q(\mem[100][1] )
         );
  EDFFX1 \mem_reg[100][0]  ( .D(n872), .E(n996), .CK(clk), .Q(\mem[100][0] )
         );
  EDFFX1 \mem_reg[104][7]  ( .D(n908), .E(n1005), .CK(clk), .Q(\mem[104][7] )
         );
  EDFFX1 \mem_reg[104][6]  ( .D(n903), .E(n1005), .CK(clk), .Q(\mem[104][6] )
         );
  EDFFX1 \mem_reg[104][5]  ( .D(n898), .E(n1005), .CK(clk), .Q(\mem[104][5] )
         );
  EDFFX1 \mem_reg[104][4]  ( .D(n893), .E(n1005), .CK(clk), .Q(\mem[104][4] )
         );
  EDFFX1 \mem_reg[104][3]  ( .D(n888), .E(n1005), .CK(clk), .Q(\mem[104][3] )
         );
  EDFFX1 \mem_reg[104][2]  ( .D(n883), .E(n1005), .CK(clk), .Q(\mem[104][2] )
         );
  EDFFX1 \mem_reg[104][1]  ( .D(n878), .E(n1005), .CK(clk), .Q(\mem[104][1] )
         );
  EDFFX1 \mem_reg[104][0]  ( .D(n873), .E(n1005), .CK(clk), .Q(\mem[104][0] )
         );
  EDFFX1 \mem_reg[108][7]  ( .D(n908), .E(n1014), .CK(clk), .Q(\mem[108][7] )
         );
  EDFFX1 \mem_reg[108][6]  ( .D(n903), .E(n1014), .CK(clk), .Q(\mem[108][6] )
         );
  EDFFX1 \mem_reg[108][5]  ( .D(n898), .E(n1014), .CK(clk), .Q(\mem[108][5] )
         );
  EDFFX1 \mem_reg[108][4]  ( .D(n893), .E(n1014), .CK(clk), .Q(\mem[108][4] )
         );
  EDFFX1 \mem_reg[108][3]  ( .D(n888), .E(n1014), .CK(clk), .Q(\mem[108][3] )
         );
  EDFFX1 \mem_reg[108][2]  ( .D(n883), .E(n1014), .CK(clk), .Q(\mem[108][2] )
         );
  EDFFX1 \mem_reg[108][1]  ( .D(n878), .E(n1014), .CK(clk), .Q(\mem[108][1] )
         );
  EDFFX1 \mem_reg[108][0]  ( .D(n873), .E(n1014), .CK(clk), .Q(\mem[108][0] )
         );
  EDFFX1 \mem_reg[112][7]  ( .D(n908), .E(n986), .CK(clk), .Q(\mem[112][7] )
         );
  EDFFX1 \mem_reg[112][6]  ( .D(n903), .E(n986), .CK(clk), .Q(\mem[112][6] )
         );
  EDFFX1 \mem_reg[112][5]  ( .D(n898), .E(n986), .CK(clk), .Q(\mem[112][5] )
         );
  EDFFX1 \mem_reg[112][4]  ( .D(n893), .E(n986), .CK(clk), .Q(\mem[112][4] )
         );
  EDFFX1 \mem_reg[112][3]  ( .D(n888), .E(n986), .CK(clk), .Q(\mem[112][3] )
         );
  EDFFX1 \mem_reg[112][2]  ( .D(n883), .E(n986), .CK(clk), .Q(\mem[112][2] )
         );
  EDFFX1 \mem_reg[112][1]  ( .D(n878), .E(n986), .CK(clk), .Q(\mem[112][1] )
         );
  EDFFX1 \mem_reg[112][0]  ( .D(n873), .E(n986), .CK(clk), .Q(\mem[112][0] )
         );
  EDFFX1 \mem_reg[116][7]  ( .D(n907), .E(n995), .CK(clk), .Q(\mem[116][7] )
         );
  EDFFX1 \mem_reg[116][6]  ( .D(n902), .E(n995), .CK(clk), .Q(\mem[116][6] )
         );
  EDFFX1 \mem_reg[116][5]  ( .D(n897), .E(n995), .CK(clk), .Q(\mem[116][5] )
         );
  EDFFX1 \mem_reg[116][4]  ( .D(n892), .E(n995), .CK(clk), .Q(\mem[116][4] )
         );
  EDFFX1 \mem_reg[116][3]  ( .D(n887), .E(n995), .CK(clk), .Q(\mem[116][3] )
         );
  EDFFX1 \mem_reg[116][2]  ( .D(n882), .E(n995), .CK(clk), .Q(\mem[116][2] )
         );
  EDFFX1 \mem_reg[116][1]  ( .D(n877), .E(n995), .CK(clk), .Q(\mem[116][1] )
         );
  EDFFX1 \mem_reg[116][0]  ( .D(n872), .E(n995), .CK(clk), .Q(\mem[116][0] )
         );
  EDFFX1 \mem_reg[120][7]  ( .D(n907), .E(n1004), .CK(clk), .Q(\mem[120][7] )
         );
  EDFFX1 \mem_reg[120][6]  ( .D(n902), .E(n1004), .CK(clk), .Q(\mem[120][6] )
         );
  EDFFX1 \mem_reg[120][5]  ( .D(n897), .E(n1004), .CK(clk), .Q(\mem[120][5] )
         );
  EDFFX1 \mem_reg[120][4]  ( .D(n892), .E(n1004), .CK(clk), .Q(\mem[120][4] )
         );
  EDFFX1 \mem_reg[120][3]  ( .D(n887), .E(n1004), .CK(clk), .Q(\mem[120][3] )
         );
  EDFFX1 \mem_reg[120][2]  ( .D(n882), .E(n1004), .CK(clk), .Q(\mem[120][2] )
         );
  EDFFX1 \mem_reg[120][1]  ( .D(n877), .E(n1004), .CK(clk), .Q(\mem[120][1] )
         );
  EDFFX1 \mem_reg[120][0]  ( .D(n872), .E(n1004), .CK(clk), .Q(\mem[120][0] )
         );
  EDFFX1 \mem_reg[124][7]  ( .D(n907), .E(n1013), .CK(clk), .Q(\mem[124][7] )
         );
  EDFFX1 \mem_reg[124][6]  ( .D(n902), .E(n1013), .CK(clk), .Q(\mem[124][6] )
         );
  EDFFX1 \mem_reg[124][5]  ( .D(n897), .E(n1013), .CK(clk), .Q(\mem[124][5] )
         );
  EDFFX1 \mem_reg[124][4]  ( .D(n892), .E(n1013), .CK(clk), .Q(\mem[124][4] )
         );
  EDFFX1 \mem_reg[124][3]  ( .D(n887), .E(n1013), .CK(clk), .Q(\mem[124][3] )
         );
  EDFFX1 \mem_reg[124][2]  ( .D(n882), .E(n1013), .CK(clk), .Q(\mem[124][2] )
         );
  EDFFX1 \mem_reg[124][1]  ( .D(n877), .E(n1013), .CK(clk), .Q(\mem[124][1] )
         );
  EDFFX1 \mem_reg[124][0]  ( .D(n872), .E(n1013), .CK(clk), .Q(\mem[124][0] )
         );
  EDFFX1 \mem_reg[2][7]  ( .D(n910), .E(n1029), .CK(clk), .Q(\mem[2][7] ) );
  EDFFX1 \mem_reg[2][6]  ( .D(n905), .E(n1029), .CK(clk), .Q(\mem[2][6] ) );
  EDFFX1 \mem_reg[2][5]  ( .D(n900), .E(n1029), .CK(clk), .Q(\mem[2][5] ) );
  EDFFX1 \mem_reg[2][4]  ( .D(n895), .E(n1029), .CK(clk), .Q(\mem[2][4] ) );
  EDFFX1 \mem_reg[2][3]  ( .D(n890), .E(n1029), .CK(clk), .Q(\mem[2][3] ) );
  EDFFX1 \mem_reg[2][2]  ( .D(n885), .E(n1029), .CK(clk), .Q(\mem[2][2] ) );
  EDFFX1 \mem_reg[2][1]  ( .D(n880), .E(n1029), .CK(clk), .Q(\mem[2][1] ) );
  EDFFX1 \mem_reg[2][0]  ( .D(n875), .E(n1029), .CK(clk), .Q(\mem[2][0] ) );
  EDFFX1 \mem_reg[6][7]  ( .D(n911), .E(n1038), .CK(clk), .Q(\mem[6][7] ) );
  EDFFX1 \mem_reg[6][6]  ( .D(n906), .E(n1038), .CK(clk), .Q(\mem[6][6] ) );
  EDFFX1 \mem_reg[6][5]  ( .D(n901), .E(n1038), .CK(clk), .Q(\mem[6][5] ) );
  EDFFX1 \mem_reg[6][4]  ( .D(n896), .E(n1038), .CK(clk), .Q(\mem[6][4] ) );
  EDFFX1 \mem_reg[6][3]  ( .D(n891), .E(n1038), .CK(clk), .Q(\mem[6][3] ) );
  EDFFX1 \mem_reg[6][2]  ( .D(n886), .E(n1038), .CK(clk), .Q(\mem[6][2] ) );
  EDFFX1 \mem_reg[6][1]  ( .D(n881), .E(n1038), .CK(clk), .Q(\mem[6][1] ) );
  EDFFX1 \mem_reg[6][0]  ( .D(n876), .E(n1038), .CK(clk), .Q(\mem[6][0] ) );
  EDFFX1 \mem_reg[10][7]  ( .D(n907), .E(n1047), .CK(clk), .Q(\mem[10][7] ) );
  EDFFX1 \mem_reg[10][6]  ( .D(n902), .E(n1047), .CK(clk), .Q(\mem[10][6] ) );
  EDFFX1 \mem_reg[10][5]  ( .D(n897), .E(n1047), .CK(clk), .Q(\mem[10][5] ) );
  EDFFX1 \mem_reg[10][4]  ( .D(n892), .E(n1047), .CK(clk), .Q(\mem[10][4] ) );
  EDFFX1 \mem_reg[10][3]  ( .D(n887), .E(n1047), .CK(clk), .Q(\mem[10][3] ) );
  EDFFX1 \mem_reg[10][2]  ( .D(n882), .E(n1047), .CK(clk), .Q(\mem[10][2] ) );
  EDFFX1 \mem_reg[10][1]  ( .D(n877), .E(n1047), .CK(clk), .Q(\mem[10][1] ) );
  EDFFX1 \mem_reg[10][0]  ( .D(n872), .E(n1047), .CK(clk), .Q(\mem[10][0] ) );
  EDFFX1 \mem_reg[14][7]  ( .D(n908), .E(n1056), .CK(clk), .Q(\mem[14][7] ) );
  EDFFX1 \mem_reg[14][6]  ( .D(n903), .E(n1056), .CK(clk), .Q(\mem[14][6] ) );
  EDFFX1 \mem_reg[14][5]  ( .D(n898), .E(n1056), .CK(clk), .Q(\mem[14][5] ) );
  EDFFX1 \mem_reg[14][4]  ( .D(n893), .E(n1056), .CK(clk), .Q(\mem[14][4] ) );
  EDFFX1 \mem_reg[14][3]  ( .D(n888), .E(n1056), .CK(clk), .Q(\mem[14][3] ) );
  EDFFX1 \mem_reg[14][2]  ( .D(n883), .E(n1056), .CK(clk), .Q(\mem[14][2] ) );
  EDFFX1 \mem_reg[14][1]  ( .D(n878), .E(n1056), .CK(clk), .Q(\mem[14][1] ) );
  EDFFX1 \mem_reg[14][0]  ( .D(n873), .E(n1056), .CK(clk), .Q(\mem[14][0] ) );
  EDFFX1 \mem_reg[18][7]  ( .D(n908), .E(n1028), .CK(clk), .Q(\mem[18][7] ) );
  EDFFX1 \mem_reg[18][6]  ( .D(n903), .E(n1028), .CK(clk), .Q(\mem[18][6] ) );
  EDFFX1 \mem_reg[18][5]  ( .D(n898), .E(n1028), .CK(clk), .Q(\mem[18][5] ) );
  EDFFX1 \mem_reg[18][4]  ( .D(n893), .E(n1028), .CK(clk), .Q(\mem[18][4] ) );
  EDFFX1 \mem_reg[18][3]  ( .D(n888), .E(n1028), .CK(clk), .Q(\mem[18][3] ) );
  EDFFX1 \mem_reg[18][2]  ( .D(n883), .E(n1028), .CK(clk), .Q(\mem[18][2] ) );
  EDFFX1 \mem_reg[18][1]  ( .D(n878), .E(n1028), .CK(clk), .Q(\mem[18][1] ) );
  EDFFX1 \mem_reg[18][0]  ( .D(n873), .E(n1028), .CK(clk), .Q(\mem[18][0] ) );
  EDFFX1 \mem_reg[22][7]  ( .D(data_in[7]), .E(n1037), .CK(clk), .Q(
        \mem[22][7] ) );
  EDFFX1 \mem_reg[22][6]  ( .D(data_in[6]), .E(n1037), .CK(clk), .Q(
        \mem[22][6] ) );
  EDFFX1 \mem_reg[22][5]  ( .D(data_in[5]), .E(n1037), .CK(clk), .Q(
        \mem[22][5] ) );
  EDFFX1 \mem_reg[22][4]  ( .D(data_in[4]), .E(n1037), .CK(clk), .Q(
        \mem[22][4] ) );
  EDFFX1 \mem_reg[22][3]  ( .D(data_in[3]), .E(n1037), .CK(clk), .Q(
        \mem[22][3] ) );
  EDFFX1 \mem_reg[22][2]  ( .D(data_in[2]), .E(n1037), .CK(clk), .Q(
        \mem[22][2] ) );
  EDFFX1 \mem_reg[22][1]  ( .D(data_in[1]), .E(n1037), .CK(clk), .Q(
        \mem[22][1] ) );
  EDFFX1 \mem_reg[22][0]  ( .D(data_in[0]), .E(n1037), .CK(clk), .Q(
        \mem[22][0] ) );
  EDFFX1 \mem_reg[26][7]  ( .D(data_in[7]), .E(n1046), .CK(clk), .Q(
        \mem[26][7] ) );
  EDFFX1 \mem_reg[26][6]  ( .D(data_in[6]), .E(n1046), .CK(clk), .Q(
        \mem[26][6] ) );
  EDFFX1 \mem_reg[26][5]  ( .D(data_in[5]), .E(n1046), .CK(clk), .Q(
        \mem[26][5] ) );
  EDFFX1 \mem_reg[26][4]  ( .D(data_in[4]), .E(n1046), .CK(clk), .Q(
        \mem[26][4] ) );
  EDFFX1 \mem_reg[26][3]  ( .D(data_in[3]), .E(n1046), .CK(clk), .Q(
        \mem[26][3] ) );
  EDFFX1 \mem_reg[26][2]  ( .D(data_in[2]), .E(n1046), .CK(clk), .Q(
        \mem[26][2] ) );
  EDFFX1 \mem_reg[26][1]  ( .D(data_in[1]), .E(n1046), .CK(clk), .Q(
        \mem[26][1] ) );
  EDFFX1 \mem_reg[26][0]  ( .D(data_in[0]), .E(n1046), .CK(clk), .Q(
        \mem[26][0] ) );
  EDFFX1 \mem_reg[30][7]  ( .D(data_in[7]), .E(n1055), .CK(clk), .Q(
        \mem[30][7] ) );
  EDFFX1 \mem_reg[30][6]  ( .D(data_in[6]), .E(n1055), .CK(clk), .Q(
        \mem[30][6] ) );
  EDFFX1 \mem_reg[30][5]  ( .D(data_in[5]), .E(n1055), .CK(clk), .Q(
        \mem[30][5] ) );
  EDFFX1 \mem_reg[30][4]  ( .D(data_in[4]), .E(n1055), .CK(clk), .Q(
        \mem[30][4] ) );
  EDFFX1 \mem_reg[30][3]  ( .D(data_in[3]), .E(n1055), .CK(clk), .Q(
        \mem[30][3] ) );
  EDFFX1 \mem_reg[30][2]  ( .D(data_in[2]), .E(n1055), .CK(clk), .Q(
        \mem[30][2] ) );
  EDFFX1 \mem_reg[30][1]  ( .D(data_in[1]), .E(n1055), .CK(clk), .Q(
        \mem[30][1] ) );
  EDFFX1 \mem_reg[30][0]  ( .D(data_in[0]), .E(n1055), .CK(clk), .Q(
        \mem[30][0] ) );
  EDFFX1 \mem_reg[34][7]  ( .D(n911), .E(n1027), .CK(clk), .Q(\mem[34][7] ) );
  EDFFX1 \mem_reg[34][6]  ( .D(n906), .E(n1027), .CK(clk), .Q(\mem[34][6] ) );
  EDFFX1 \mem_reg[34][5]  ( .D(n901), .E(n1027), .CK(clk), .Q(\mem[34][5] ) );
  EDFFX1 \mem_reg[34][4]  ( .D(n896), .E(n1027), .CK(clk), .Q(\mem[34][4] ) );
  EDFFX1 \mem_reg[34][3]  ( .D(n891), .E(n1027), .CK(clk), .Q(\mem[34][3] ) );
  EDFFX1 \mem_reg[34][2]  ( .D(n886), .E(n1027), .CK(clk), .Q(\mem[34][2] ) );
  EDFFX1 \mem_reg[34][1]  ( .D(n881), .E(n1027), .CK(clk), .Q(\mem[34][1] ) );
  EDFFX1 \mem_reg[34][0]  ( .D(n876), .E(n1027), .CK(clk), .Q(\mem[34][0] ) );
  EDFFX1 \mem_reg[38][7]  ( .D(n911), .E(n1036), .CK(clk), .Q(\mem[38][7] ) );
  EDFFX1 \mem_reg[38][6]  ( .D(n906), .E(n1036), .CK(clk), .Q(\mem[38][6] ) );
  EDFFX1 \mem_reg[38][5]  ( .D(n901), .E(n1036), .CK(clk), .Q(\mem[38][5] ) );
  EDFFX1 \mem_reg[38][4]  ( .D(n896), .E(n1036), .CK(clk), .Q(\mem[38][4] ) );
  EDFFX1 \mem_reg[38][3]  ( .D(n891), .E(n1036), .CK(clk), .Q(\mem[38][3] ) );
  EDFFX1 \mem_reg[38][2]  ( .D(n886), .E(n1036), .CK(clk), .Q(\mem[38][2] ) );
  EDFFX1 \mem_reg[38][1]  ( .D(n881), .E(n1036), .CK(clk), .Q(\mem[38][1] ) );
  EDFFX1 \mem_reg[38][0]  ( .D(n876), .E(n1036), .CK(clk), .Q(\mem[38][0] ) );
  EDFFX1 \mem_reg[42][7]  ( .D(n911), .E(n1045), .CK(clk), .Q(\mem[42][7] ) );
  EDFFX1 \mem_reg[42][6]  ( .D(n906), .E(n1045), .CK(clk), .Q(\mem[42][6] ) );
  EDFFX1 \mem_reg[42][5]  ( .D(n901), .E(n1045), .CK(clk), .Q(\mem[42][5] ) );
  EDFFX1 \mem_reg[42][4]  ( .D(n896), .E(n1045), .CK(clk), .Q(\mem[42][4] ) );
  EDFFX1 \mem_reg[42][3]  ( .D(n891), .E(n1045), .CK(clk), .Q(\mem[42][3] ) );
  EDFFX1 \mem_reg[42][2]  ( .D(n886), .E(n1045), .CK(clk), .Q(\mem[42][2] ) );
  EDFFX1 \mem_reg[42][1]  ( .D(n881), .E(n1045), .CK(clk), .Q(\mem[42][1] ) );
  EDFFX1 \mem_reg[42][0]  ( .D(n876), .E(n1045), .CK(clk), .Q(\mem[42][0] ) );
  EDFFX1 \mem_reg[46][7]  ( .D(n908), .E(n1054), .CK(clk), .Q(\mem[46][7] ) );
  EDFFX1 \mem_reg[46][6]  ( .D(n903), .E(n1054), .CK(clk), .Q(\mem[46][6] ) );
  EDFFX1 \mem_reg[46][5]  ( .D(n898), .E(n1054), .CK(clk), .Q(\mem[46][5] ) );
  EDFFX1 \mem_reg[46][4]  ( .D(n893), .E(n1054), .CK(clk), .Q(\mem[46][4] ) );
  EDFFX1 \mem_reg[46][3]  ( .D(n888), .E(n1054), .CK(clk), .Q(\mem[46][3] ) );
  EDFFX1 \mem_reg[46][2]  ( .D(n883), .E(n1054), .CK(clk), .Q(\mem[46][2] ) );
  EDFFX1 \mem_reg[46][1]  ( .D(n878), .E(n1054), .CK(clk), .Q(\mem[46][1] ) );
  EDFFX1 \mem_reg[46][0]  ( .D(n873), .E(n1054), .CK(clk), .Q(\mem[46][0] ) );
  EDFFX1 \mem_reg[50][7]  ( .D(n908), .E(n1026), .CK(clk), .Q(\mem[50][7] ) );
  EDFFX1 \mem_reg[50][6]  ( .D(n903), .E(n1026), .CK(clk), .Q(\mem[50][6] ) );
  EDFFX1 \mem_reg[50][5]  ( .D(n898), .E(n1026), .CK(clk), .Q(\mem[50][5] ) );
  EDFFX1 \mem_reg[50][4]  ( .D(n893), .E(n1026), .CK(clk), .Q(\mem[50][4] ) );
  EDFFX1 \mem_reg[50][3]  ( .D(n888), .E(n1026), .CK(clk), .Q(\mem[50][3] ) );
  EDFFX1 \mem_reg[50][2]  ( .D(n883), .E(n1026), .CK(clk), .Q(\mem[50][2] ) );
  EDFFX1 \mem_reg[50][1]  ( .D(n878), .E(n1026), .CK(clk), .Q(\mem[50][1] ) );
  EDFFX1 \mem_reg[50][0]  ( .D(n873), .E(n1026), .CK(clk), .Q(\mem[50][0] ) );
  EDFFX1 \mem_reg[54][7]  ( .D(n911), .E(n1035), .CK(clk), .Q(\mem[54][7] ) );
  EDFFX1 \mem_reg[54][6]  ( .D(n906), .E(n1035), .CK(clk), .Q(\mem[54][6] ) );
  EDFFX1 \mem_reg[54][5]  ( .D(n901), .E(n1035), .CK(clk), .Q(\mem[54][5] ) );
  EDFFX1 \mem_reg[54][4]  ( .D(n896), .E(n1035), .CK(clk), .Q(\mem[54][4] ) );
  EDFFX1 \mem_reg[54][3]  ( .D(n891), .E(n1035), .CK(clk), .Q(\mem[54][3] ) );
  EDFFX1 \mem_reg[54][2]  ( .D(n886), .E(n1035), .CK(clk), .Q(\mem[54][2] ) );
  EDFFX1 \mem_reg[54][1]  ( .D(n881), .E(n1035), .CK(clk), .Q(\mem[54][1] ) );
  EDFFX1 \mem_reg[54][0]  ( .D(n876), .E(n1035), .CK(clk), .Q(\mem[54][0] ) );
  EDFFX1 \mem_reg[58][7]  ( .D(n910), .E(n1044), .CK(clk), .Q(\mem[58][7] ) );
  EDFFX1 \mem_reg[58][6]  ( .D(n905), .E(n1044), .CK(clk), .Q(\mem[58][6] ) );
  EDFFX1 \mem_reg[58][5]  ( .D(n900), .E(n1044), .CK(clk), .Q(\mem[58][5] ) );
  EDFFX1 \mem_reg[58][4]  ( .D(n895), .E(n1044), .CK(clk), .Q(\mem[58][4] ) );
  EDFFX1 \mem_reg[58][3]  ( .D(n890), .E(n1044), .CK(clk), .Q(\mem[58][3] ) );
  EDFFX1 \mem_reg[58][2]  ( .D(n885), .E(n1044), .CK(clk), .Q(\mem[58][2] ) );
  EDFFX1 \mem_reg[58][1]  ( .D(n880), .E(n1044), .CK(clk), .Q(\mem[58][1] ) );
  EDFFX1 \mem_reg[58][0]  ( .D(n875), .E(n1044), .CK(clk), .Q(\mem[58][0] ) );
  EDFFX1 \mem_reg[62][7]  ( .D(n910), .E(n1053), .CK(clk), .Q(\mem[62][7] ) );
  EDFFX1 \mem_reg[62][6]  ( .D(n905), .E(n1053), .CK(clk), .Q(\mem[62][6] ) );
  EDFFX1 \mem_reg[62][5]  ( .D(n900), .E(n1053), .CK(clk), .Q(\mem[62][5] ) );
  EDFFX1 \mem_reg[62][4]  ( .D(n895), .E(n1053), .CK(clk), .Q(\mem[62][4] ) );
  EDFFX1 \mem_reg[62][3]  ( .D(n890), .E(n1053), .CK(clk), .Q(\mem[62][3] ) );
  EDFFX1 \mem_reg[62][2]  ( .D(n885), .E(n1053), .CK(clk), .Q(\mem[62][2] ) );
  EDFFX1 \mem_reg[62][1]  ( .D(n880), .E(n1053), .CK(clk), .Q(\mem[62][1] ) );
  EDFFX1 \mem_reg[62][0]  ( .D(n875), .E(n1053), .CK(clk), .Q(\mem[62][0] ) );
  EDFFX1 \mem_reg[66][7]  ( .D(n910), .E(n1025), .CK(clk), .Q(\mem[66][7] ) );
  EDFFX1 \mem_reg[66][6]  ( .D(n905), .E(n1025), .CK(clk), .Q(\mem[66][6] ) );
  EDFFX1 \mem_reg[66][5]  ( .D(n900), .E(n1025), .CK(clk), .Q(\mem[66][5] ) );
  EDFFX1 \mem_reg[66][4]  ( .D(n895), .E(n1025), .CK(clk), .Q(\mem[66][4] ) );
  EDFFX1 \mem_reg[66][3]  ( .D(n890), .E(n1025), .CK(clk), .Q(\mem[66][3] ) );
  EDFFX1 \mem_reg[66][2]  ( .D(n885), .E(n1025), .CK(clk), .Q(\mem[66][2] ) );
  EDFFX1 \mem_reg[66][1]  ( .D(n880), .E(n1025), .CK(clk), .Q(\mem[66][1] ) );
  EDFFX1 \mem_reg[66][0]  ( .D(n875), .E(n1025), .CK(clk), .Q(\mem[66][0] ) );
  EDFFX1 \mem_reg[70][7]  ( .D(n909), .E(n1034), .CK(clk), .Q(\mem[70][7] ) );
  EDFFX1 \mem_reg[70][6]  ( .D(n904), .E(n1034), .CK(clk), .Q(\mem[70][6] ) );
  EDFFX1 \mem_reg[70][5]  ( .D(n899), .E(n1034), .CK(clk), .Q(\mem[70][5] ) );
  EDFFX1 \mem_reg[70][4]  ( .D(n894), .E(n1034), .CK(clk), .Q(\mem[70][4] ) );
  EDFFX1 \mem_reg[70][3]  ( .D(n889), .E(n1034), .CK(clk), .Q(\mem[70][3] ) );
  EDFFX1 \mem_reg[70][2]  ( .D(n884), .E(n1034), .CK(clk), .Q(\mem[70][2] ) );
  EDFFX1 \mem_reg[70][1]  ( .D(n879), .E(n1034), .CK(clk), .Q(\mem[70][1] ) );
  EDFFX1 \mem_reg[70][0]  ( .D(n874), .E(n1034), .CK(clk), .Q(\mem[70][0] ) );
  EDFFX1 \mem_reg[74][7]  ( .D(n909), .E(n1043), .CK(clk), .Q(\mem[74][7] ) );
  EDFFX1 \mem_reg[74][6]  ( .D(n904), .E(n1043), .CK(clk), .Q(\mem[74][6] ) );
  EDFFX1 \mem_reg[74][5]  ( .D(n899), .E(n1043), .CK(clk), .Q(\mem[74][5] ) );
  EDFFX1 \mem_reg[74][4]  ( .D(n894), .E(n1043), .CK(clk), .Q(\mem[74][4] ) );
  EDFFX1 \mem_reg[74][3]  ( .D(n889), .E(n1043), .CK(clk), .Q(\mem[74][3] ) );
  EDFFX1 \mem_reg[74][2]  ( .D(n884), .E(n1043), .CK(clk), .Q(\mem[74][2] ) );
  EDFFX1 \mem_reg[74][1]  ( .D(n879), .E(n1043), .CK(clk), .Q(\mem[74][1] ) );
  EDFFX1 \mem_reg[74][0]  ( .D(n874), .E(n1043), .CK(clk), .Q(\mem[74][0] ) );
  EDFFX1 \mem_reg[78][7]  ( .D(n909), .E(n1052), .CK(clk), .Q(\mem[78][7] ) );
  EDFFX1 \mem_reg[78][6]  ( .D(n904), .E(n1052), .CK(clk), .Q(\mem[78][6] ) );
  EDFFX1 \mem_reg[78][5]  ( .D(n899), .E(n1052), .CK(clk), .Q(\mem[78][5] ) );
  EDFFX1 \mem_reg[78][4]  ( .D(n894), .E(n1052), .CK(clk), .Q(\mem[78][4] ) );
  EDFFX1 \mem_reg[78][3]  ( .D(n889), .E(n1052), .CK(clk), .Q(\mem[78][3] ) );
  EDFFX1 \mem_reg[78][2]  ( .D(n884), .E(n1052), .CK(clk), .Q(\mem[78][2] ) );
  EDFFX1 \mem_reg[78][1]  ( .D(n879), .E(n1052), .CK(clk), .Q(\mem[78][1] ) );
  EDFFX1 \mem_reg[78][0]  ( .D(n874), .E(n1052), .CK(clk), .Q(\mem[78][0] ) );
  EDFFX1 \mem_reg[82][7]  ( .D(n909), .E(n1024), .CK(clk), .Q(\mem[82][7] ) );
  EDFFX1 \mem_reg[82][6]  ( .D(n904), .E(n1024), .CK(clk), .Q(\mem[82][6] ) );
  EDFFX1 \mem_reg[82][5]  ( .D(n899), .E(n1024), .CK(clk), .Q(\mem[82][5] ) );
  EDFFX1 \mem_reg[82][4]  ( .D(n894), .E(n1024), .CK(clk), .Q(\mem[82][4] ) );
  EDFFX1 \mem_reg[82][3]  ( .D(n889), .E(n1024), .CK(clk), .Q(\mem[82][3] ) );
  EDFFX1 \mem_reg[82][2]  ( .D(n884), .E(n1024), .CK(clk), .Q(\mem[82][2] ) );
  EDFFX1 \mem_reg[82][1]  ( .D(n879), .E(n1024), .CK(clk), .Q(\mem[82][1] ) );
  EDFFX1 \mem_reg[82][0]  ( .D(n874), .E(n1024), .CK(clk), .Q(\mem[82][0] ) );
  EDFFX1 \mem_reg[86][7]  ( .D(n909), .E(n1033), .CK(clk), .Q(\mem[86][7] ) );
  EDFFX1 \mem_reg[86][6]  ( .D(n904), .E(n1033), .CK(clk), .Q(\mem[86][6] ) );
  EDFFX1 \mem_reg[86][5]  ( .D(n899), .E(n1033), .CK(clk), .Q(\mem[86][5] ) );
  EDFFX1 \mem_reg[86][4]  ( .D(n894), .E(n1033), .CK(clk), .Q(\mem[86][4] ) );
  EDFFX1 \mem_reg[86][3]  ( .D(n889), .E(n1033), .CK(clk), .Q(\mem[86][3] ) );
  EDFFX1 \mem_reg[86][2]  ( .D(n884), .E(n1033), .CK(clk), .Q(\mem[86][2] ) );
  EDFFX1 \mem_reg[86][1]  ( .D(n879), .E(n1033), .CK(clk), .Q(\mem[86][1] ) );
  EDFFX1 \mem_reg[86][0]  ( .D(n874), .E(n1033), .CK(clk), .Q(\mem[86][0] ) );
  EDFFX1 \mem_reg[90][7]  ( .D(n909), .E(n1042), .CK(clk), .Q(\mem[90][7] ) );
  EDFFX1 \mem_reg[90][6]  ( .D(n904), .E(n1042), .CK(clk), .Q(\mem[90][6] ) );
  EDFFX1 \mem_reg[90][5]  ( .D(n899), .E(n1042), .CK(clk), .Q(\mem[90][5] ) );
  EDFFX1 \mem_reg[90][4]  ( .D(n894), .E(n1042), .CK(clk), .Q(\mem[90][4] ) );
  EDFFX1 \mem_reg[90][3]  ( .D(n889), .E(n1042), .CK(clk), .Q(\mem[90][3] ) );
  EDFFX1 \mem_reg[90][2]  ( .D(n884), .E(n1042), .CK(clk), .Q(\mem[90][2] ) );
  EDFFX1 \mem_reg[90][1]  ( .D(n879), .E(n1042), .CK(clk), .Q(\mem[90][1] ) );
  EDFFX1 \mem_reg[90][0]  ( .D(n874), .E(n1042), .CK(clk), .Q(\mem[90][0] ) );
  EDFFX1 \mem_reg[94][7]  ( .D(n908), .E(n1051), .CK(clk), .Q(\mem[94][7] ) );
  EDFFX1 \mem_reg[94][6]  ( .D(n903), .E(n1051), .CK(clk), .Q(\mem[94][6] ) );
  EDFFX1 \mem_reg[94][5]  ( .D(n898), .E(n1051), .CK(clk), .Q(\mem[94][5] ) );
  EDFFX1 \mem_reg[94][4]  ( .D(n893), .E(n1051), .CK(clk), .Q(\mem[94][4] ) );
  EDFFX1 \mem_reg[94][3]  ( .D(n888), .E(n1051), .CK(clk), .Q(\mem[94][3] ) );
  EDFFX1 \mem_reg[94][2]  ( .D(n883), .E(n1051), .CK(clk), .Q(\mem[94][2] ) );
  EDFFX1 \mem_reg[94][1]  ( .D(n878), .E(n1051), .CK(clk), .Q(\mem[94][1] ) );
  EDFFX1 \mem_reg[94][0]  ( .D(n873), .E(n1051), .CK(clk), .Q(\mem[94][0] ) );
  EDFFX1 \mem_reg[98][7]  ( .D(n910), .E(n1023), .CK(clk), .Q(\mem[98][7] ) );
  EDFFX1 \mem_reg[98][6]  ( .D(n905), .E(n1023), .CK(clk), .Q(\mem[98][6] ) );
  EDFFX1 \mem_reg[98][5]  ( .D(n900), .E(n1023), .CK(clk), .Q(\mem[98][5] ) );
  EDFFX1 \mem_reg[98][4]  ( .D(n895), .E(n1023), .CK(clk), .Q(\mem[98][4] ) );
  EDFFX1 \mem_reg[98][3]  ( .D(n890), .E(n1023), .CK(clk), .Q(\mem[98][3] ) );
  EDFFX1 \mem_reg[98][2]  ( .D(n885), .E(n1023), .CK(clk), .Q(\mem[98][2] ) );
  EDFFX1 \mem_reg[98][1]  ( .D(n880), .E(n1023), .CK(clk), .Q(\mem[98][1] ) );
  EDFFX1 \mem_reg[98][0]  ( .D(n875), .E(n1023), .CK(clk), .Q(\mem[98][0] ) );
  EDFFX1 \mem_reg[102][7]  ( .D(n911), .E(n1032), .CK(clk), .Q(\mem[102][7] )
         );
  EDFFX1 \mem_reg[102][6]  ( .D(n906), .E(n1032), .CK(clk), .Q(\mem[102][6] )
         );
  EDFFX1 \mem_reg[102][5]  ( .D(n901), .E(n1032), .CK(clk), .Q(\mem[102][5] )
         );
  EDFFX1 \mem_reg[102][4]  ( .D(n896), .E(n1032), .CK(clk), .Q(\mem[102][4] )
         );
  EDFFX1 \mem_reg[102][3]  ( .D(n891), .E(n1032), .CK(clk), .Q(\mem[102][3] )
         );
  EDFFX1 \mem_reg[102][2]  ( .D(n886), .E(n1032), .CK(clk), .Q(\mem[102][2] )
         );
  EDFFX1 \mem_reg[102][1]  ( .D(n881), .E(n1032), .CK(clk), .Q(\mem[102][1] )
         );
  EDFFX1 \mem_reg[102][0]  ( .D(n876), .E(n1032), .CK(clk), .Q(\mem[102][0] )
         );
  EDFFX1 \mem_reg[106][7]  ( .D(n908), .E(n1041), .CK(clk), .Q(\mem[106][7] )
         );
  EDFFX1 \mem_reg[106][6]  ( .D(n903), .E(n1041), .CK(clk), .Q(\mem[106][6] )
         );
  EDFFX1 \mem_reg[106][5]  ( .D(n898), .E(n1041), .CK(clk), .Q(\mem[106][5] )
         );
  EDFFX1 \mem_reg[106][4]  ( .D(n893), .E(n1041), .CK(clk), .Q(\mem[106][4] )
         );
  EDFFX1 \mem_reg[106][3]  ( .D(n888), .E(n1041), .CK(clk), .Q(\mem[106][3] )
         );
  EDFFX1 \mem_reg[106][2]  ( .D(n883), .E(n1041), .CK(clk), .Q(\mem[106][2] )
         );
  EDFFX1 \mem_reg[106][1]  ( .D(n878), .E(n1041), .CK(clk), .Q(\mem[106][1] )
         );
  EDFFX1 \mem_reg[106][0]  ( .D(n873), .E(n1041), .CK(clk), .Q(\mem[106][0] )
         );
  EDFFX1 \mem_reg[110][7]  ( .D(n908), .E(n1050), .CK(clk), .Q(\mem[110][7] )
         );
  EDFFX1 \mem_reg[110][6]  ( .D(n903), .E(n1050), .CK(clk), .Q(\mem[110][6] )
         );
  EDFFX1 \mem_reg[110][5]  ( .D(n898), .E(n1050), .CK(clk), .Q(\mem[110][5] )
         );
  EDFFX1 \mem_reg[110][4]  ( .D(n893), .E(n1050), .CK(clk), .Q(\mem[110][4] )
         );
  EDFFX1 \mem_reg[110][3]  ( .D(n888), .E(n1050), .CK(clk), .Q(\mem[110][3] )
         );
  EDFFX1 \mem_reg[110][2]  ( .D(n883), .E(n1050), .CK(clk), .Q(\mem[110][2] )
         );
  EDFFX1 \mem_reg[110][1]  ( .D(n878), .E(n1050), .CK(clk), .Q(\mem[110][1] )
         );
  EDFFX1 \mem_reg[110][0]  ( .D(n873), .E(n1050), .CK(clk), .Q(\mem[110][0] )
         );
  EDFFX1 \mem_reg[114][7]  ( .D(n908), .E(n1022), .CK(clk), .Q(\mem[114][7] )
         );
  EDFFX1 \mem_reg[114][6]  ( .D(n903), .E(n1022), .CK(clk), .Q(\mem[114][6] )
         );
  EDFFX1 \mem_reg[114][5]  ( .D(n898), .E(n1022), .CK(clk), .Q(\mem[114][5] )
         );
  EDFFX1 \mem_reg[114][4]  ( .D(n893), .E(n1022), .CK(clk), .Q(\mem[114][4] )
         );
  EDFFX1 \mem_reg[114][3]  ( .D(n888), .E(n1022), .CK(clk), .Q(\mem[114][3] )
         );
  EDFFX1 \mem_reg[114][2]  ( .D(n883), .E(n1022), .CK(clk), .Q(\mem[114][2] )
         );
  EDFFX1 \mem_reg[114][1]  ( .D(n878), .E(n1022), .CK(clk), .Q(\mem[114][1] )
         );
  EDFFX1 \mem_reg[114][0]  ( .D(n873), .E(n1022), .CK(clk), .Q(\mem[114][0] )
         );
  EDFFX1 \mem_reg[118][7]  ( .D(n907), .E(n1031), .CK(clk), .Q(\mem[118][7] )
         );
  EDFFX1 \mem_reg[118][6]  ( .D(n902), .E(n1031), .CK(clk), .Q(\mem[118][6] )
         );
  EDFFX1 \mem_reg[118][5]  ( .D(n897), .E(n1031), .CK(clk), .Q(\mem[118][5] )
         );
  EDFFX1 \mem_reg[118][4]  ( .D(n892), .E(n1031), .CK(clk), .Q(\mem[118][4] )
         );
  EDFFX1 \mem_reg[118][3]  ( .D(n887), .E(n1031), .CK(clk), .Q(\mem[118][3] )
         );
  EDFFX1 \mem_reg[118][2]  ( .D(n882), .E(n1031), .CK(clk), .Q(\mem[118][2] )
         );
  EDFFX1 \mem_reg[118][1]  ( .D(n877), .E(n1031), .CK(clk), .Q(\mem[118][1] )
         );
  EDFFX1 \mem_reg[118][0]  ( .D(n872), .E(n1031), .CK(clk), .Q(\mem[118][0] )
         );
  EDFFX1 \mem_reg[122][7]  ( .D(n907), .E(n1040), .CK(clk), .Q(\mem[122][7] )
         );
  EDFFX1 \mem_reg[122][6]  ( .D(n902), .E(n1040), .CK(clk), .Q(\mem[122][6] )
         );
  EDFFX1 \mem_reg[122][5]  ( .D(n897), .E(n1040), .CK(clk), .Q(\mem[122][5] )
         );
  EDFFX1 \mem_reg[122][4]  ( .D(n892), .E(n1040), .CK(clk), .Q(\mem[122][4] )
         );
  EDFFX1 \mem_reg[122][3]  ( .D(n887), .E(n1040), .CK(clk), .Q(\mem[122][3] )
         );
  EDFFX1 \mem_reg[122][2]  ( .D(n882), .E(n1040), .CK(clk), .Q(\mem[122][2] )
         );
  EDFFX1 \mem_reg[122][1]  ( .D(n877), .E(n1040), .CK(clk), .Q(\mem[122][1] )
         );
  EDFFX1 \mem_reg[122][0]  ( .D(n872), .E(n1040), .CK(clk), .Q(\mem[122][0] )
         );
  EDFFX1 \mem_reg[126][7]  ( .D(n907), .E(n1049), .CK(clk), .Q(\mem[126][7] )
         );
  EDFFX1 \mem_reg[126][6]  ( .D(n902), .E(n1049), .CK(clk), .Q(\mem[126][6] )
         );
  EDFFX1 \mem_reg[126][5]  ( .D(n897), .E(n1049), .CK(clk), .Q(\mem[126][5] )
         );
  EDFFX1 \mem_reg[126][4]  ( .D(n892), .E(n1049), .CK(clk), .Q(\mem[126][4] )
         );
  EDFFX1 \mem_reg[126][3]  ( .D(n887), .E(n1049), .CK(clk), .Q(\mem[126][3] )
         );
  EDFFX1 \mem_reg[126][2]  ( .D(n882), .E(n1049), .CK(clk), .Q(\mem[126][2] )
         );
  EDFFX1 \mem_reg[126][1]  ( .D(n877), .E(n1049), .CK(clk), .Q(\mem[126][1] )
         );
  EDFFX1 \mem_reg[126][0]  ( .D(n872), .E(n1049), .CK(clk), .Q(\mem[126][0] )
         );
  DFFRX1 \valid_mem_reg[127]  ( .D(n448), .CK(clk), .RN(n3), .Q(valid_mem[127]) );
  DFFRX1 \valid_mem_reg[111]  ( .D(n464), .CK(clk), .RN(n4), .Q(valid_mem[111]) );
  DFFRX1 \valid_mem_reg[110]  ( .D(n465), .CK(clk), .RN(n3), .Q(valid_mem[110]) );
  DFFRX1 \valid_mem_reg[109]  ( .D(n466), .CK(clk), .RN(n4), .Q(valid_mem[109]) );
  DFFRX1 \valid_mem_reg[108]  ( .D(n467), .CK(clk), .RN(n3), .Q(valid_mem[108]) );
  DFFRX1 \valid_mem_reg[107]  ( .D(n468), .CK(clk), .RN(n4), .Q(valid_mem[107]) );
  DFFRX1 \valid_mem_reg[106]  ( .D(n469), .CK(clk), .RN(n3), .Q(valid_mem[106]) );
  DFFRX1 \valid_mem_reg[105]  ( .D(n470), .CK(clk), .RN(n4), .Q(valid_mem[105]) );
  DFFRX1 \valid_mem_reg[104]  ( .D(n471), .CK(clk), .RN(n3), .Q(valid_mem[104]) );
  DFFRX1 \valid_mem_reg[103]  ( .D(n472), .CK(clk), .RN(n4), .Q(valid_mem[103]) );
  DFFRX1 \valid_mem_reg[102]  ( .D(n473), .CK(clk), .RN(n3), .Q(valid_mem[102]) );
  DFFRX1 \valid_mem_reg[101]  ( .D(n474), .CK(clk), .RN(n4), .Q(valid_mem[101]) );
  DFFRX1 \valid_mem_reg[100]  ( .D(n475), .CK(clk), .RN(n3), .Q(valid_mem[100]) );
  DFFRX1 \valid_mem_reg[99]  ( .D(n476), .CK(clk), .RN(n4), .Q(valid_mem[99])
         );
  DFFRX1 \valid_mem_reg[98]  ( .D(n477), .CK(clk), .RN(n3), .Q(valid_mem[98])
         );
  DFFRX1 \valid_mem_reg[97]  ( .D(n478), .CK(clk), .RN(n4), .Q(valid_mem[97])
         );
  DFFRX1 \valid_mem_reg[96]  ( .D(n479), .CK(clk), .RN(n3), .Q(valid_mem[96])
         );
  DFFRX1 \valid_mem_reg[95]  ( .D(n480), .CK(clk), .RN(n4), .Q(valid_mem[95])
         );
  DFFRX1 \valid_mem_reg[94]  ( .D(n481), .CK(clk), .RN(n3), .Q(valid_mem[94])
         );
  DFFRX1 \valid_mem_reg[93]  ( .D(n482), .CK(clk), .RN(n4), .Q(valid_mem[93])
         );
  DFFRX1 \valid_mem_reg[92]  ( .D(n483), .CK(clk), .RN(n3), .Q(valid_mem[92])
         );
  DFFRX1 \valid_mem_reg[91]  ( .D(n484), .CK(clk), .RN(n4), .Q(valid_mem[91])
         );
  DFFRX1 \valid_mem_reg[90]  ( .D(n485), .CK(clk), .RN(n3), .Q(valid_mem[90])
         );
  DFFRX1 \valid_mem_reg[89]  ( .D(n486), .CK(clk), .RN(n4), .Q(valid_mem[89])
         );
  DFFRX1 \valid_mem_reg[88]  ( .D(n487), .CK(clk), .RN(n3), .Q(valid_mem[88])
         );
  DFFRX1 \valid_mem_reg[87]  ( .D(n488), .CK(clk), .RN(n4), .Q(valid_mem[87])
         );
  DFFRX1 \valid_mem_reg[86]  ( .D(n489), .CK(clk), .RN(n3), .Q(valid_mem[86])
         );
  DFFRX1 \valid_mem_reg[85]  ( .D(n490), .CK(clk), .RN(n4), .Q(valid_mem[85])
         );
  DFFRX1 \valid_mem_reg[84]  ( .D(n491), .CK(clk), .RN(n3), .Q(valid_mem[84])
         );
  DFFRX1 \valid_mem_reg[83]  ( .D(n492), .CK(clk), .RN(n4), .Q(valid_mem[83])
         );
  DFFRX1 \valid_mem_reg[82]  ( .D(n493), .CK(clk), .RN(n3), .Q(valid_mem[82])
         );
  DFFRX1 \valid_mem_reg[81]  ( .D(n494), .CK(clk), .RN(n4), .Q(valid_mem[81])
         );
  DFFRX1 \valid_mem_reg[80]  ( .D(n495), .CK(clk), .RN(n3), .Q(valid_mem[80])
         );
  DFFRX1 \valid_mem_reg[79]  ( .D(n496), .CK(clk), .RN(n4), .Q(valid_mem[79])
         );
  DFFRX1 \valid_mem_reg[78]  ( .D(n497), .CK(clk), .RN(n3), .Q(valid_mem[78])
         );
  DFFRX1 \valid_mem_reg[77]  ( .D(n498), .CK(clk), .RN(n4), .Q(valid_mem[77])
         );
  DFFRX1 \valid_mem_reg[76]  ( .D(n499), .CK(clk), .RN(n3), .Q(valid_mem[76])
         );
  DFFRX1 \valid_mem_reg[75]  ( .D(n500), .CK(clk), .RN(n4), .Q(valid_mem[75])
         );
  DFFRX1 \valid_mem_reg[74]  ( .D(n501), .CK(clk), .RN(n3), .Q(valid_mem[74])
         );
  DFFRX1 \valid_mem_reg[73]  ( .D(n502), .CK(clk), .RN(n4), .Q(valid_mem[73])
         );
  DFFRX1 \valid_mem_reg[72]  ( .D(n503), .CK(clk), .RN(n3), .Q(valid_mem[72])
         );
  DFFRX1 \valid_mem_reg[71]  ( .D(n504), .CK(clk), .RN(n4), .Q(valid_mem[71])
         );
  DFFRX1 \valid_mem_reg[70]  ( .D(n505), .CK(clk), .RN(n3), .Q(valid_mem[70])
         );
  DFFRX1 \valid_mem_reg[69]  ( .D(n506), .CK(clk), .RN(n4), .Q(valid_mem[69])
         );
  DFFRX1 \valid_mem_reg[68]  ( .D(n507), .CK(clk), .RN(n3), .Q(valid_mem[68])
         );
  DFFRX1 \valid_mem_reg[67]  ( .D(n508), .CK(clk), .RN(n4), .Q(valid_mem[67])
         );
  DFFRX1 \valid_mem_reg[66]  ( .D(n509), .CK(clk), .RN(n3), .Q(valid_mem[66])
         );
  DFFRX1 \valid_mem_reg[65]  ( .D(n510), .CK(clk), .RN(n4), .Q(valid_mem[65])
         );
  DFFRX1 \valid_mem_reg[64]  ( .D(n511), .CK(clk), .RN(n3), .Q(valid_mem[64])
         );
  DFFRX1 \valid_mem_reg[63]  ( .D(n512), .CK(clk), .RN(n4), .Q(valid_mem[63])
         );
  DFFRX1 \valid_mem_reg[62]  ( .D(n513), .CK(clk), .RN(n3), .Q(valid_mem[62])
         );
  DFFRX1 \valid_mem_reg[61]  ( .D(n514), .CK(clk), .RN(n4), .Q(valid_mem[61])
         );
  DFFRX1 \valid_mem_reg[60]  ( .D(n515), .CK(clk), .RN(n3), .Q(valid_mem[60])
         );
  DFFRX1 \valid_mem_reg[59]  ( .D(n516), .CK(clk), .RN(n4), .Q(valid_mem[59])
         );
  DFFRX1 \valid_mem_reg[58]  ( .D(n517), .CK(clk), .RN(n3), .Q(valid_mem[58])
         );
  DFFRX1 \valid_mem_reg[57]  ( .D(n518), .CK(clk), .RN(n4), .Q(valid_mem[57])
         );
  DFFRX1 \valid_mem_reg[56]  ( .D(n519), .CK(clk), .RN(n3), .Q(valid_mem[56])
         );
  DFFRX1 \valid_mem_reg[55]  ( .D(n520), .CK(clk), .RN(n4), .Q(valid_mem[55])
         );
  DFFRX1 \valid_mem_reg[54]  ( .D(n521), .CK(clk), .RN(n3), .Q(valid_mem[54])
         );
  DFFRX1 \valid_mem_reg[53]  ( .D(n522), .CK(clk), .RN(n4), .Q(valid_mem[53])
         );
  DFFRX1 \valid_mem_reg[52]  ( .D(n523), .CK(clk), .RN(n3), .Q(valid_mem[52])
         );
  DFFRX1 \valid_mem_reg[51]  ( .D(n524), .CK(clk), .RN(n4), .Q(valid_mem[51])
         );
  DFFRX1 \valid_mem_reg[50]  ( .D(n525), .CK(clk), .RN(n3), .Q(valid_mem[50])
         );
  DFFRX1 \valid_mem_reg[49]  ( .D(n526), .CK(clk), .RN(n4), .Q(valid_mem[49])
         );
  DFFRX1 \valid_mem_reg[48]  ( .D(n527), .CK(clk), .RN(n3), .Q(valid_mem[48])
         );
  DFFRX1 \valid_mem_reg[47]  ( .D(n528), .CK(clk), .RN(n4), .Q(valid_mem[47])
         );
  DFFRX1 \valid_mem_reg[46]  ( .D(n529), .CK(clk), .RN(n3), .Q(valid_mem[46])
         );
  DFFRX1 \valid_mem_reg[45]  ( .D(n530), .CK(clk), .RN(n4), .Q(valid_mem[45])
         );
  DFFRX1 \valid_mem_reg[44]  ( .D(n531), .CK(clk), .RN(n3), .Q(valid_mem[44])
         );
  DFFRX1 \valid_mem_reg[43]  ( .D(n532), .CK(clk), .RN(n4), .Q(valid_mem[43])
         );
  DFFRX1 \valid_mem_reg[42]  ( .D(n533), .CK(clk), .RN(n3), .Q(valid_mem[42])
         );
  DFFRX1 \valid_mem_reg[41]  ( .D(n534), .CK(clk), .RN(n4), .Q(valid_mem[41])
         );
  DFFRX1 \valid_mem_reg[40]  ( .D(n535), .CK(clk), .RN(n3), .Q(valid_mem[40])
         );
  DFFRX1 \valid_mem_reg[39]  ( .D(n536), .CK(clk), .RN(n4), .Q(valid_mem[39])
         );
  DFFRX1 \valid_mem_reg[38]  ( .D(n537), .CK(clk), .RN(n3), .Q(valid_mem[38])
         );
  DFFRX1 \valid_mem_reg[37]  ( .D(n538), .CK(clk), .RN(n4), .Q(valid_mem[37])
         );
  DFFRX1 \valid_mem_reg[36]  ( .D(n539), .CK(clk), .RN(n3), .Q(valid_mem[36])
         );
  DFFRX1 \valid_mem_reg[35]  ( .D(n540), .CK(clk), .RN(n4), .Q(valid_mem[35])
         );
  DFFRX1 \valid_mem_reg[34]  ( .D(n541), .CK(clk), .RN(n3), .Q(valid_mem[34])
         );
  DFFRX1 \valid_mem_reg[33]  ( .D(n542), .CK(clk), .RN(n4), .Q(valid_mem[33])
         );
  DFFRX1 \valid_mem_reg[32]  ( .D(n543), .CK(clk), .RN(n3), .Q(valid_mem[32])
         );
  DFFRX1 \valid_mem_reg[31]  ( .D(n544), .CK(clk), .RN(n4), .Q(valid_mem[31])
         );
  DFFRX1 \valid_mem_reg[30]  ( .D(n545), .CK(clk), .RN(n3), .Q(valid_mem[30])
         );
  DFFRX1 \valid_mem_reg[29]  ( .D(n546), .CK(clk), .RN(n4), .Q(valid_mem[29])
         );
  DFFRX1 \valid_mem_reg[28]  ( .D(n547), .CK(clk), .RN(n3), .Q(valid_mem[28])
         );
  DFFRX1 \valid_mem_reg[27]  ( .D(n548), .CK(clk), .RN(n4), .Q(valid_mem[27])
         );
  DFFRX1 \valid_mem_reg[26]  ( .D(n549), .CK(clk), .RN(n3), .Q(valid_mem[26])
         );
  DFFRX1 \valid_mem_reg[25]  ( .D(n550), .CK(clk), .RN(n4), .Q(valid_mem[25])
         );
  DFFRX1 \valid_mem_reg[24]  ( .D(n551), .CK(clk), .RN(n3), .Q(valid_mem[24])
         );
  DFFRX1 \valid_mem_reg[23]  ( .D(n552), .CK(clk), .RN(n4), .Q(valid_mem[23])
         );
  DFFRX1 \valid_mem_reg[22]  ( .D(n553), .CK(clk), .RN(n3), .Q(valid_mem[22])
         );
  DFFRX1 \valid_mem_reg[21]  ( .D(n554), .CK(clk), .RN(n4), .Q(valid_mem[21])
         );
  DFFRX1 \valid_mem_reg[20]  ( .D(n555), .CK(clk), .RN(n3), .Q(valid_mem[20])
         );
  DFFRX1 \valid_mem_reg[19]  ( .D(n556), .CK(clk), .RN(n4), .Q(valid_mem[19])
         );
  DFFRX1 \valid_mem_reg[18]  ( .D(n557), .CK(clk), .RN(n3), .Q(valid_mem[18])
         );
  DFFRX1 \valid_mem_reg[17]  ( .D(n558), .CK(clk), .RN(n4), .Q(valid_mem[17])
         );
  DFFRX1 \valid_mem_reg[16]  ( .D(n559), .CK(clk), .RN(n3), .Q(valid_mem[16])
         );
  DFFRX1 \valid_mem_reg[15]  ( .D(n560), .CK(clk), .RN(n4), .Q(valid_mem[15])
         );
  DFFRX1 \valid_mem_reg[14]  ( .D(n561), .CK(clk), .RN(n3), .Q(valid_mem[14])
         );
  DFFRX1 \valid_mem_reg[13]  ( .D(n562), .CK(clk), .RN(n4), .Q(valid_mem[13])
         );
  DFFRX1 \valid_mem_reg[12]  ( .D(n563), .CK(clk), .RN(n3), .Q(valid_mem[12])
         );
  DFFRX1 \valid_mem_reg[11]  ( .D(n564), .CK(clk), .RN(n4), .Q(valid_mem[11])
         );
  DFFRX1 \valid_mem_reg[10]  ( .D(n565), .CK(clk), .RN(n3), .Q(valid_mem[10])
         );
  DFFRX1 \valid_mem_reg[9]  ( .D(n566), .CK(clk), .RN(n4), .Q(valid_mem[9]) );
  DFFRX1 \valid_mem_reg[8]  ( .D(n567), .CK(clk), .RN(n3), .Q(valid_mem[8]) );
  DFFRX1 \valid_mem_reg[7]  ( .D(n568), .CK(clk), .RN(n4), .Q(valid_mem[7]) );
  DFFRX1 \valid_mem_reg[6]  ( .D(n569), .CK(clk), .RN(n3), .Q(valid_mem[6]) );
  DFFRX1 \valid_mem_reg[5]  ( .D(n570), .CK(clk), .RN(n4), .Q(valid_mem[5]) );
  DFFRX1 \valid_mem_reg[4]  ( .D(n571), .CK(clk), .RN(n3), .Q(valid_mem[4]) );
  DFFRX1 \valid_mem_reg[3]  ( .D(n572), .CK(clk), .RN(n4), .Q(valid_mem[3]) );
  DFFRX1 \valid_mem_reg[2]  ( .D(n573), .CK(clk), .RN(n3), .Q(valid_mem[2]) );
  DFFRX1 \valid_mem_reg[1]  ( .D(n574), .CK(clk), .RN(n4), .Q(valid_mem[1]) );
  DFFRX1 \valid_mem_reg[0]  ( .D(n575), .CK(clk), .RN(n3), .Q(valid_mem[0]) );
  DFFRX1 \valid_mem_reg[126]  ( .D(n449), .CK(clk), .RN(n4), .Q(valid_mem[126]) );
  DFFRX1 \valid_mem_reg[125]  ( .D(n450), .CK(clk), .RN(n3), .Q(valid_mem[125]) );
  DFFRX1 \valid_mem_reg[124]  ( .D(n451), .CK(clk), .RN(n4), .Q(valid_mem[124]) );
  DFFRX1 \valid_mem_reg[123]  ( .D(n452), .CK(clk), .RN(n3), .Q(valid_mem[123]) );
  DFFRX1 \valid_mem_reg[122]  ( .D(n453), .CK(clk), .RN(n4), .Q(valid_mem[122]) );
  DFFRX1 \valid_mem_reg[121]  ( .D(n454), .CK(clk), .RN(n3), .Q(valid_mem[121]) );
  DFFRX1 \valid_mem_reg[120]  ( .D(n455), .CK(clk), .RN(n4), .Q(valid_mem[120]) );
  DFFRX1 \valid_mem_reg[119]  ( .D(n456), .CK(clk), .RN(n3), .Q(valid_mem[119]) );
  DFFRX1 \valid_mem_reg[118]  ( .D(n457), .CK(clk), .RN(n4), .Q(valid_mem[118]) );
  DFFRX1 \valid_mem_reg[117]  ( .D(n458), .CK(clk), .RN(n3), .Q(valid_mem[117]) );
  DFFRX1 \valid_mem_reg[116]  ( .D(n459), .CK(clk), .RN(n4), .Q(valid_mem[116]) );
  DFFRX1 \valid_mem_reg[115]  ( .D(n460), .CK(clk), .RN(n3), .Q(valid_mem[115]) );
  DFFRX1 \valid_mem_reg[114]  ( .D(n461), .CK(clk), .RN(n4), .Q(valid_mem[114]) );
  DFFRX1 \valid_mem_reg[113]  ( .D(n462), .CK(clk), .RN(n3), .Q(valid_mem[113]) );
  DFFRX1 \valid_mem_reg[112]  ( .D(n463), .CK(clk), .RN(n4), .Q(valid_mem[112]) );
  DFFRX1 valid_reg ( .D(N41), .CK(clk), .RN(n3), .QN(n1) );
  DFFRX1 \data_out_reg[7]  ( .D(N33), .CK(clk), .RN(n4), .Q(data_out[7]) );
  DFFRX1 \data_out_reg[6]  ( .D(N34), .CK(clk), .RN(n3), .Q(data_out[6]) );
  DFFRX1 \data_out_reg[5]  ( .D(N35), .CK(clk), .RN(n4), .Q(data_out[5]) );
  DFFRX1 \data_out_reg[4]  ( .D(N36), .CK(clk), .RN(n3), .Q(data_out[4]) );
  DFFRX1 \data_out_reg[3]  ( .D(N37), .CK(clk), .RN(n4), .Q(data_out[3]) );
  DFFRX1 \data_out_reg[2]  ( .D(N38), .CK(clk), .RN(n3), .Q(data_out[2]) );
  DFFRX1 \data_out_reg[1]  ( .D(N39), .CK(clk), .RN(n4), .Q(data_out[1]) );
  DFFRX1 \data_out_reg[0]  ( .D(N40), .CK(clk), .RN(n3), .Q(data_out[0]) );
  NOR2BX4 U3 ( .AN(n912), .B(n269), .Y(n865) );
  NOR2BX4 U4 ( .AN(n912), .B(n302), .Y(n863) );
  NOR2BX4 U5 ( .AN(n912), .B(n335), .Y(n861) );
  NOR2BX4 U6 ( .AN(n912), .B(n368), .Y(n859) );
  NOR2BX4 U7 ( .AN(n912), .B(n401), .Y(n857) );
  INVX4 U8 ( .A(n1), .Y(valid) );
  INVX12 U9 ( .A(rst), .Y(n3) );
  INVX12 U10 ( .A(rst), .Y(n4) );
  CLKBUFX3 U11 ( .A(n433), .Y(n869) );
  CLKBUFX3 U12 ( .A(n434), .Y(n867) );
  CLKBUFX3 U13 ( .A(n432), .Y(n871) );
  NOR2X1 U14 ( .A(n1058), .B(n985), .Y(n441) );
  NOR2X1 U15 ( .A(n1060), .B(n1059), .Y(n440) );
  NOR2X1 U16 ( .A(n1058), .B(write_counter_count[0]), .Y(n442) );
  NOR2X1 U17 ( .A(n1059), .B(write_counter_count[3]), .Y(n446) );
  NOR2X1 U18 ( .A(n1060), .B(write_counter_count[2]), .Y(n445) );
  NOR2X1 U19 ( .A(n985), .B(write_counter_count[1]), .Y(n443) );
  NOR2X1 U20 ( .A(write_counter_count[0]), .B(write_counter_count[1]), .Y(n444) );
  NOR2X1 U21 ( .A(write_counter_count[2]), .B(write_counter_count[3]), .Y(n447) );
  CLKBUFX3 U22 ( .A(n828), .Y(n840) );
  CLKBUFX3 U23 ( .A(n827), .Y(n842) );
  CLKBUFX3 U24 ( .A(n828), .Y(n841) );
  CLKBUFX3 U25 ( .A(n828), .Y(n839) );
  CLKBUFX3 U26 ( .A(n830), .Y(n838) );
  CLKBUFX3 U27 ( .A(n830), .Y(n837) );
  CLKBUFX3 U28 ( .A(n829), .Y(n836) );
  CLKBUFX3 U29 ( .A(n829), .Y(n835) );
  CLKBUFX3 U30 ( .A(n830), .Y(n833) );
  CLKBUFX3 U31 ( .A(n830), .Y(n834) );
  CLKBUFX3 U32 ( .A(n830), .Y(n831) );
  CLKBUFX3 U33 ( .A(n829), .Y(n832) );
  CLKBUFX3 U34 ( .A(n803), .Y(n825) );
  CLKBUFX3 U35 ( .A(n803), .Y(n824) );
  CLKBUFX3 U36 ( .A(n803), .Y(n821) );
  CLKBUFX3 U37 ( .A(n804), .Y(n823) );
  CLKBUFX3 U38 ( .A(n803), .Y(n822) );
  CLKBUFX3 U39 ( .A(n803), .Y(n819) );
  CLKBUFX3 U40 ( .A(n803), .Y(n820) );
  CLKBUFX3 U41 ( .A(n804), .Y(n816) );
  CLKBUFX3 U42 ( .A(n803), .Y(n818) );
  CLKBUFX3 U43 ( .A(n804), .Y(n817) );
  CLKBUFX3 U44 ( .A(n802), .Y(n814) );
  CLKBUFX3 U45 ( .A(n804), .Y(n815) );
  CLKBUFX3 U46 ( .A(n803), .Y(n811) );
  CLKBUFX3 U47 ( .A(n805), .Y(n813) );
  CLKBUFX3 U48 ( .A(n804), .Y(n812) );
  CLKBUFX3 U49 ( .A(n804), .Y(n809) );
  CLKBUFX3 U50 ( .A(n804), .Y(n810) );
  CLKBUFX3 U51 ( .A(n805), .Y(n806) );
  CLKBUFX3 U52 ( .A(n803), .Y(n807) );
  CLKBUFX3 U53 ( .A(n804), .Y(n808) );
  CLKBUFX3 U54 ( .A(n827), .Y(n843) );
  CLKBUFX3 U55 ( .A(n826), .Y(n827) );
  CLKBUFX3 U56 ( .A(n826), .Y(n828) );
  CLKBUFX3 U57 ( .A(N27), .Y(n829) );
  CLKBUFX3 U58 ( .A(n826), .Y(n830) );
  INVX3 U59 ( .A(n152), .Y(n940) );
  INVX3 U60 ( .A(n201), .Y(n941) );
  INVX3 U61 ( .A(n204), .Y(n1050) );
  INVX3 U62 ( .A(n206), .Y(n977) );
  INVX3 U63 ( .A(n208), .Y(n1014) );
  INVX3 U64 ( .A(n210), .Y(n932) );
  INVX3 U65 ( .A(n212), .Y(n1041) );
  INVX3 U66 ( .A(n214), .Y(n968) );
  INVX3 U67 ( .A(n216), .Y(n1005) );
  INVX3 U68 ( .A(n218), .Y(n923) );
  INVX3 U69 ( .A(n220), .Y(n1032) );
  INVX3 U70 ( .A(n222), .Y(n959) );
  INVX3 U71 ( .A(n224), .Y(n996) );
  INVX3 U72 ( .A(n226), .Y(n914) );
  INVX3 U73 ( .A(n228), .Y(n1023) );
  INVX3 U74 ( .A(n230), .Y(n950) );
  INVX3 U75 ( .A(n232), .Y(n987) );
  INVX3 U76 ( .A(n234), .Y(n942) );
  INVX3 U77 ( .A(n237), .Y(n1051) );
  INVX3 U78 ( .A(n239), .Y(n978) );
  INVX3 U79 ( .A(n241), .Y(n1015) );
  INVX3 U80 ( .A(n243), .Y(n933) );
  INVX3 U81 ( .A(n245), .Y(n1042) );
  INVX3 U82 ( .A(n247), .Y(n969) );
  INVX3 U83 ( .A(n249), .Y(n1006) );
  INVX3 U84 ( .A(n251), .Y(n924) );
  INVX3 U85 ( .A(n253), .Y(n1033) );
  INVX3 U86 ( .A(n255), .Y(n960) );
  INVX3 U87 ( .A(n257), .Y(n997) );
  INVX3 U88 ( .A(n259), .Y(n915) );
  INVX3 U89 ( .A(n261), .Y(n1024) );
  INVX3 U90 ( .A(n263), .Y(n951) );
  INVX3 U91 ( .A(n265), .Y(n988) );
  INVX3 U92 ( .A(n267), .Y(n943) );
  INVX3 U93 ( .A(n270), .Y(n1052) );
  INVX3 U94 ( .A(n272), .Y(n979) );
  INVX3 U95 ( .A(n274), .Y(n1016) );
  INVX3 U96 ( .A(n276), .Y(n934) );
  INVX3 U97 ( .A(n278), .Y(n1043) );
  INVX3 U98 ( .A(n280), .Y(n970) );
  INVX3 U99 ( .A(n282), .Y(n1007) );
  INVX3 U100 ( .A(n284), .Y(n925) );
  INVX3 U101 ( .A(n286), .Y(n1034) );
  INVX3 U102 ( .A(n288), .Y(n961) );
  INVX3 U103 ( .A(n290), .Y(n998) );
  INVX3 U104 ( .A(n292), .Y(n916) );
  INVX3 U105 ( .A(n294), .Y(n1025) );
  INVX3 U106 ( .A(n296), .Y(n952) );
  INVX3 U107 ( .A(n298), .Y(n989) );
  INVX3 U108 ( .A(n300), .Y(n944) );
  INVX3 U109 ( .A(n303), .Y(n1053) );
  INVX3 U110 ( .A(n305), .Y(n980) );
  INVX3 U111 ( .A(n307), .Y(n1017) );
  INVX3 U112 ( .A(n309), .Y(n935) );
  INVX3 U113 ( .A(n311), .Y(n1044) );
  INVX3 U114 ( .A(n313), .Y(n971) );
  INVX3 U115 ( .A(n315), .Y(n1008) );
  INVX3 U116 ( .A(n317), .Y(n926) );
  INVX3 U117 ( .A(n319), .Y(n1035) );
  INVX3 U118 ( .A(n321), .Y(n962) );
  INVX3 U119 ( .A(n323), .Y(n999) );
  INVX3 U120 ( .A(n325), .Y(n917) );
  INVX3 U121 ( .A(n327), .Y(n1026) );
  INVX3 U122 ( .A(n329), .Y(n953) );
  INVX3 U123 ( .A(n331), .Y(n990) );
  INVX3 U124 ( .A(n333), .Y(n945) );
  INVX3 U125 ( .A(n336), .Y(n1054) );
  INVX3 U126 ( .A(n338), .Y(n981) );
  INVX3 U127 ( .A(n340), .Y(n1018) );
  INVX3 U128 ( .A(n342), .Y(n936) );
  INVX3 U129 ( .A(n344), .Y(n1045) );
  INVX3 U130 ( .A(n346), .Y(n972) );
  INVX3 U131 ( .A(n348), .Y(n1009) );
  INVX3 U132 ( .A(n350), .Y(n927) );
  INVX3 U133 ( .A(n352), .Y(n1036) );
  INVX3 U134 ( .A(n354), .Y(n963) );
  INVX3 U135 ( .A(n356), .Y(n1000) );
  INVX3 U136 ( .A(n358), .Y(n918) );
  INVX3 U137 ( .A(n360), .Y(n1027) );
  INVX3 U138 ( .A(n362), .Y(n954) );
  INVX3 U139 ( .A(n364), .Y(n991) );
  INVX3 U140 ( .A(n366), .Y(n946) );
  INVX3 U141 ( .A(n369), .Y(n1055) );
  INVX3 U142 ( .A(n371), .Y(n982) );
  INVX3 U143 ( .A(n373), .Y(n1019) );
  INVX3 U144 ( .A(n375), .Y(n937) );
  INVX3 U145 ( .A(n377), .Y(n1046) );
  INVX3 U146 ( .A(n379), .Y(n973) );
  INVX3 U147 ( .A(n381), .Y(n1010) );
  INVX3 U148 ( .A(n383), .Y(n928) );
  INVX3 U149 ( .A(n385), .Y(n1037) );
  INVX3 U150 ( .A(n387), .Y(n964) );
  INVX3 U151 ( .A(n389), .Y(n1001) );
  INVX3 U152 ( .A(n391), .Y(n919) );
  INVX3 U153 ( .A(n393), .Y(n1028) );
  INVX3 U154 ( .A(n395), .Y(n955) );
  INVX3 U155 ( .A(n397), .Y(n992) );
  INVX3 U156 ( .A(n399), .Y(n947) );
  INVX3 U157 ( .A(n402), .Y(n1056) );
  INVX3 U158 ( .A(n404), .Y(n983) );
  INVX3 U159 ( .A(n406), .Y(n1020) );
  INVX3 U160 ( .A(n408), .Y(n938) );
  INVX3 U161 ( .A(n410), .Y(n1047) );
  INVX3 U162 ( .A(n412), .Y(n974) );
  INVX3 U163 ( .A(n414), .Y(n1011) );
  INVX3 U164 ( .A(n416), .Y(n929) );
  INVX3 U165 ( .A(n418), .Y(n1038) );
  INVX3 U166 ( .A(n420), .Y(n965) );
  INVX3 U167 ( .A(n422), .Y(n1002) );
  INVX3 U168 ( .A(n424), .Y(n920) );
  INVX3 U169 ( .A(n426), .Y(n1029) );
  INVX3 U170 ( .A(n428), .Y(n956) );
  INVX3 U171 ( .A(n430), .Y(n993) );
  INVX3 U172 ( .A(n156), .Y(n1049) );
  INVX3 U173 ( .A(n159), .Y(n976) );
  INVX3 U174 ( .A(n162), .Y(n1013) );
  INVX3 U175 ( .A(n165), .Y(n931) );
  INVX3 U176 ( .A(n168), .Y(n1040) );
  INVX3 U177 ( .A(n171), .Y(n967) );
  INVX3 U178 ( .A(n174), .Y(n1004) );
  INVX3 U179 ( .A(n177), .Y(n922) );
  INVX3 U180 ( .A(n180), .Y(n1031) );
  INVX3 U181 ( .A(n183), .Y(n958) );
  INVX3 U182 ( .A(n186), .Y(n995) );
  INVX3 U183 ( .A(n189), .Y(n913) );
  INVX3 U184 ( .A(n192), .Y(n1022) );
  INVX3 U185 ( .A(n195), .Y(n949) );
  INVX3 U186 ( .A(n198), .Y(n986) );
  INVX3 U187 ( .A(n155), .Y(n948) );
  CLKBUFX3 U188 ( .A(n848), .Y(n852) );
  CLKBUFX3 U189 ( .A(n848), .Y(n851) );
  CLKBUFX3 U190 ( .A(n848), .Y(n850) );
  CLKBUFX3 U191 ( .A(n848), .Y(n849) );
  CLKBUFX3 U192 ( .A(n844), .Y(n847) );
  CLKBUFX3 U193 ( .A(n844), .Y(n846) );
  CLKBUFX3 U194 ( .A(n844), .Y(n845) );
  CLKBUFX3 U195 ( .A(data_in[0]), .Y(n873) );
  CLKBUFX3 U196 ( .A(data_in[1]), .Y(n878) );
  CLKBUFX3 U197 ( .A(data_in[2]), .Y(n883) );
  CLKBUFX3 U198 ( .A(data_in[3]), .Y(n888) );
  CLKBUFX3 U199 ( .A(data_in[4]), .Y(n893) );
  CLKBUFX3 U200 ( .A(data_in[5]), .Y(n898) );
  CLKBUFX3 U201 ( .A(data_in[6]), .Y(n903) );
  CLKBUFX3 U202 ( .A(data_in[7]), .Y(n908) );
  CLKBUFX3 U203 ( .A(data_in[0]), .Y(n874) );
  CLKBUFX3 U204 ( .A(data_in[1]), .Y(n879) );
  CLKBUFX3 U205 ( .A(data_in[2]), .Y(n884) );
  CLKBUFX3 U206 ( .A(data_in[3]), .Y(n889) );
  CLKBUFX3 U207 ( .A(data_in[4]), .Y(n894) );
  CLKBUFX3 U208 ( .A(data_in[5]), .Y(n899) );
  CLKBUFX3 U209 ( .A(data_in[6]), .Y(n904) );
  CLKBUFX3 U210 ( .A(data_in[7]), .Y(n909) );
  CLKBUFX3 U211 ( .A(data_in[0]), .Y(n875) );
  CLKBUFX3 U212 ( .A(data_in[1]), .Y(n880) );
  CLKBUFX3 U213 ( .A(data_in[2]), .Y(n885) );
  CLKBUFX3 U214 ( .A(data_in[3]), .Y(n890) );
  CLKBUFX3 U215 ( .A(data_in[4]), .Y(n895) );
  CLKBUFX3 U216 ( .A(data_in[5]), .Y(n900) );
  CLKBUFX3 U217 ( .A(data_in[6]), .Y(n905) );
  CLKBUFX3 U218 ( .A(data_in[7]), .Y(n910) );
  CLKBUFX3 U219 ( .A(data_in[0]), .Y(n876) );
  CLKBUFX3 U220 ( .A(data_in[1]), .Y(n881) );
  CLKBUFX3 U221 ( .A(data_in[2]), .Y(n886) );
  CLKBUFX3 U222 ( .A(data_in[3]), .Y(n891) );
  CLKBUFX3 U223 ( .A(data_in[4]), .Y(n896) );
  CLKBUFX3 U224 ( .A(data_in[5]), .Y(n901) );
  CLKBUFX3 U225 ( .A(data_in[6]), .Y(n906) );
  CLKBUFX3 U226 ( .A(data_in[7]), .Y(n911) );
  CLKBUFX3 U227 ( .A(n802), .Y(n805) );
  CLKBUFX3 U228 ( .A(N27), .Y(n826) );
  NAND2X1 U229 ( .A(n869), .B(n1057), .Y(n204) );
  NAND2X1 U230 ( .A(n869), .B(n984), .Y(n206) );
  NAND2X1 U231 ( .A(n869), .B(n1021), .Y(n208) );
  NAND2X1 U232 ( .A(n869), .B(n939), .Y(n210) );
  NAND2X1 U233 ( .A(n869), .B(n1048), .Y(n212) );
  NAND2X1 U234 ( .A(n869), .B(n975), .Y(n214) );
  NAND2X1 U235 ( .A(n869), .B(n1012), .Y(n216) );
  NAND2X1 U236 ( .A(n869), .B(n930), .Y(n218) );
  NAND2X1 U237 ( .A(n869), .B(n1039), .Y(n220) );
  NAND2X1 U238 ( .A(n869), .B(n966), .Y(n222) );
  NAND2X1 U239 ( .A(n869), .B(n1003), .Y(n224) );
  NAND2X1 U240 ( .A(n869), .B(n921), .Y(n226) );
  NAND2X1 U241 ( .A(n869), .B(n1030), .Y(n228) );
  NAND2X1 U242 ( .A(n869), .B(n957), .Y(n230) );
  NAND2X1 U243 ( .A(n869), .B(n994), .Y(n232) );
  NAND2X1 U244 ( .A(n867), .B(n1057), .Y(n237) );
  NAND2X1 U245 ( .A(n867), .B(n984), .Y(n239) );
  NAND2X1 U246 ( .A(n867), .B(n1021), .Y(n241) );
  NAND2X1 U247 ( .A(n867), .B(n939), .Y(n243) );
  NAND2X1 U248 ( .A(n867), .B(n1048), .Y(n245) );
  NAND2X1 U249 ( .A(n867), .B(n975), .Y(n247) );
  NAND2X1 U250 ( .A(n867), .B(n1012), .Y(n249) );
  NAND2X1 U251 ( .A(n867), .B(n930), .Y(n251) );
  NAND2X1 U252 ( .A(n867), .B(n1039), .Y(n253) );
  NAND2X1 U253 ( .A(n867), .B(n966), .Y(n255) );
  NAND2X1 U254 ( .A(n867), .B(n1003), .Y(n257) );
  NAND2X1 U255 ( .A(n867), .B(n921), .Y(n259) );
  NAND2X1 U256 ( .A(n867), .B(n1030), .Y(n261) );
  NAND2X1 U257 ( .A(n867), .B(n957), .Y(n263) );
  NAND2X1 U258 ( .A(n867), .B(n994), .Y(n265) );
  NAND2X1 U259 ( .A(n865), .B(n1057), .Y(n270) );
  NAND2X1 U260 ( .A(n865), .B(n984), .Y(n272) );
  NAND2X1 U261 ( .A(n865), .B(n1021), .Y(n274) );
  NAND2X1 U262 ( .A(n865), .B(n939), .Y(n276) );
  NAND2X1 U263 ( .A(n865), .B(n1048), .Y(n278) );
  NAND2X1 U264 ( .A(n865), .B(n975), .Y(n280) );
  NAND2X1 U265 ( .A(n865), .B(n1012), .Y(n282) );
  NAND2X1 U266 ( .A(n865), .B(n930), .Y(n284) );
  NAND2X1 U267 ( .A(n865), .B(n1039), .Y(n286) );
  NAND2X1 U268 ( .A(n865), .B(n966), .Y(n288) );
  NAND2X1 U269 ( .A(n865), .B(n1003), .Y(n290) );
  NAND2X1 U270 ( .A(n865), .B(n921), .Y(n292) );
  NAND2X1 U271 ( .A(n865), .B(n1030), .Y(n294) );
  NAND2X1 U272 ( .A(n865), .B(n957), .Y(n296) );
  NAND2X1 U273 ( .A(n865), .B(n994), .Y(n298) );
  NAND2X1 U274 ( .A(n863), .B(n1057), .Y(n303) );
  NAND2X1 U275 ( .A(n863), .B(n984), .Y(n305) );
  NAND2X1 U276 ( .A(n863), .B(n1021), .Y(n307) );
  NAND2X1 U277 ( .A(n863), .B(n939), .Y(n309) );
  NAND2X1 U278 ( .A(n863), .B(n1048), .Y(n311) );
  NAND2X1 U279 ( .A(n863), .B(n975), .Y(n313) );
  NAND2X1 U280 ( .A(n863), .B(n1012), .Y(n315) );
  NAND2X1 U281 ( .A(n863), .B(n930), .Y(n317) );
  NAND2X1 U282 ( .A(n863), .B(n1039), .Y(n319) );
  NAND2X1 U283 ( .A(n863), .B(n966), .Y(n321) );
  NAND2X1 U284 ( .A(n863), .B(n1003), .Y(n323) );
  NAND2X1 U285 ( .A(n863), .B(n921), .Y(n325) );
  NAND2X1 U286 ( .A(n863), .B(n1030), .Y(n327) );
  NAND2X1 U287 ( .A(n863), .B(n957), .Y(n329) );
  NAND2X1 U288 ( .A(n863), .B(n994), .Y(n331) );
  NAND2X1 U289 ( .A(n861), .B(n1057), .Y(n336) );
  NAND2X1 U290 ( .A(n861), .B(n984), .Y(n338) );
  NAND2X1 U291 ( .A(n861), .B(n1021), .Y(n340) );
  NAND2X1 U292 ( .A(n861), .B(n939), .Y(n342) );
  NAND2X1 U293 ( .A(n861), .B(n1048), .Y(n344) );
  NAND2X1 U294 ( .A(n861), .B(n975), .Y(n346) );
  NAND2X1 U295 ( .A(n861), .B(n1012), .Y(n348) );
  NAND2X1 U296 ( .A(n861), .B(n930), .Y(n350) );
  NAND2X1 U297 ( .A(n861), .B(n1039), .Y(n352) );
  NAND2X1 U298 ( .A(n861), .B(n966), .Y(n354) );
  NAND2X1 U299 ( .A(n861), .B(n1003), .Y(n356) );
  NAND2X1 U300 ( .A(n861), .B(n921), .Y(n358) );
  NAND2X1 U301 ( .A(n861), .B(n1030), .Y(n360) );
  NAND2X1 U302 ( .A(n861), .B(n957), .Y(n362) );
  NAND2X1 U303 ( .A(n861), .B(n994), .Y(n364) );
  NAND2X1 U304 ( .A(n859), .B(n1057), .Y(n369) );
  NAND2X1 U305 ( .A(n859), .B(n984), .Y(n371) );
  NAND2X1 U306 ( .A(n859), .B(n1021), .Y(n373) );
  NAND2X1 U307 ( .A(n859), .B(n939), .Y(n375) );
  NAND2X1 U308 ( .A(n859), .B(n1048), .Y(n377) );
  NAND2X1 U309 ( .A(n859), .B(n975), .Y(n379) );
  NAND2X1 U310 ( .A(n859), .B(n1012), .Y(n381) );
  NAND2X1 U311 ( .A(n859), .B(n930), .Y(n383) );
  NAND2X1 U312 ( .A(n859), .B(n1039), .Y(n385) );
  NAND2X1 U313 ( .A(n859), .B(n966), .Y(n387) );
  NAND2X1 U314 ( .A(n859), .B(n1003), .Y(n389) );
  NAND2X1 U315 ( .A(n859), .B(n921), .Y(n391) );
  NAND2X1 U316 ( .A(n859), .B(n1030), .Y(n393) );
  NAND2X1 U317 ( .A(n859), .B(n957), .Y(n395) );
  NAND2X1 U318 ( .A(n859), .B(n994), .Y(n397) );
  NAND2X1 U319 ( .A(n857), .B(n1057), .Y(n402) );
  NAND2X1 U320 ( .A(n857), .B(n984), .Y(n404) );
  NAND2X1 U321 ( .A(n857), .B(n1021), .Y(n406) );
  NAND2X1 U322 ( .A(n857), .B(n939), .Y(n408) );
  NAND2X1 U323 ( .A(n857), .B(n1048), .Y(n410) );
  NAND2X1 U324 ( .A(n857), .B(n975), .Y(n412) );
  NAND2X1 U325 ( .A(n857), .B(n1012), .Y(n414) );
  NAND2X1 U326 ( .A(n857), .B(n930), .Y(n416) );
  NAND2X1 U327 ( .A(n857), .B(n1039), .Y(n418) );
  NAND2X1 U328 ( .A(n857), .B(n966), .Y(n420) );
  NAND2X1 U329 ( .A(n857), .B(n1003), .Y(n422) );
  NAND2X1 U330 ( .A(n857), .B(n921), .Y(n424) );
  NAND2X1 U331 ( .A(n857), .B(n1030), .Y(n426) );
  NAND2X1 U332 ( .A(n857), .B(n957), .Y(n428) );
  NAND2X1 U333 ( .A(n857), .B(n994), .Y(n430) );
  NAND2X1 U334 ( .A(n871), .B(n948), .Y(n152) );
  NAND2X1 U335 ( .A(n869), .B(n948), .Y(n201) );
  NAND2X1 U336 ( .A(n867), .B(n948), .Y(n234) );
  NAND2X1 U337 ( .A(n865), .B(n948), .Y(n267) );
  NAND2X1 U338 ( .A(n863), .B(n948), .Y(n300) );
  NAND2X1 U339 ( .A(n861), .B(n948), .Y(n333) );
  NAND2X1 U340 ( .A(n859), .B(n948), .Y(n366) );
  NAND2X1 U341 ( .A(n857), .B(n948), .Y(n399) );
  NAND2X1 U342 ( .A(n1057), .B(n871), .Y(n156) );
  NAND2X1 U343 ( .A(n984), .B(n871), .Y(n159) );
  NAND2X1 U344 ( .A(n1021), .B(n871), .Y(n162) );
  NAND2X1 U345 ( .A(n939), .B(n871), .Y(n165) );
  NAND2X1 U346 ( .A(n1048), .B(n871), .Y(n168) );
  NAND2X1 U347 ( .A(n975), .B(n871), .Y(n171) );
  NAND2X1 U348 ( .A(n1012), .B(n871), .Y(n174) );
  NAND2X1 U349 ( .A(n930), .B(n871), .Y(n177) );
  NAND2X1 U350 ( .A(n1039), .B(n871), .Y(n180) );
  NAND2X1 U351 ( .A(n966), .B(n871), .Y(n183) );
  NAND2X1 U352 ( .A(n1003), .B(n871), .Y(n186) );
  NAND2X1 U353 ( .A(n921), .B(n871), .Y(n189) );
  NAND2X1 U354 ( .A(n1030), .B(n871), .Y(n192) );
  NAND2X1 U355 ( .A(n957), .B(n871), .Y(n195) );
  NAND2X1 U356 ( .A(n994), .B(n871), .Y(n198) );
  CLKBUFX3 U357 ( .A(en), .Y(n912) );
  INVX3 U358 ( .A(n170), .Y(n1048) );
  INVX3 U359 ( .A(n158), .Y(n1057) );
  INVX3 U360 ( .A(n161), .Y(n984) );
  INVX3 U361 ( .A(n164), .Y(n1021) );
  INVX3 U362 ( .A(n173), .Y(n975) );
  INVX3 U363 ( .A(n176), .Y(n1012) );
  INVX3 U364 ( .A(n182), .Y(n1039) );
  INVX3 U365 ( .A(n194), .Y(n1030) );
  INVX3 U366 ( .A(n167), .Y(n939) );
  INVX3 U367 ( .A(n179), .Y(n930) );
  INVX3 U368 ( .A(n185), .Y(n966) );
  INVX3 U369 ( .A(n188), .Y(n1003) );
  INVX3 U370 ( .A(n191), .Y(n921) );
  INVX3 U371 ( .A(n197), .Y(n957) );
  INVX3 U372 ( .A(n200), .Y(n994) );
  NAND2X2 U373 ( .A(n440), .B(n441), .Y(n155) );
  CLKBUFX3 U374 ( .A(data_in[0]), .Y(n872) );
  CLKBUFX3 U375 ( .A(data_in[1]), .Y(n877) );
  CLKBUFX3 U376 ( .A(data_in[2]), .Y(n882) );
  CLKBUFX3 U377 ( .A(data_in[3]), .Y(n887) );
  CLKBUFX3 U378 ( .A(data_in[4]), .Y(n892) );
  CLKBUFX3 U379 ( .A(data_in[5]), .Y(n897) );
  CLKBUFX3 U380 ( .A(data_in[6]), .Y(n902) );
  CLKBUFX3 U381 ( .A(data_in[7]), .Y(n907) );
  CLKBUFX3 U382 ( .A(N29), .Y(n848) );
  CLKBUFX3 U383 ( .A(N28), .Y(n844) );
  CLKBUFX3 U384 ( .A(N26), .Y(n804) );
  CLKBUFX3 U385 ( .A(N26), .Y(n803) );
  CLKBUFX3 U386 ( .A(N26), .Y(n802) );
  NOR2BX1 U387 ( .AN(n912), .B(n868), .Y(n433) );
  NOR2BX1 U388 ( .AN(n912), .B(n866), .Y(n434) );
  NOR2BX1 U389 ( .AN(n912), .B(n870), .Y(n432) );
  NAND2X2 U390 ( .A(n445), .B(n442), .Y(n170) );
  NAND2X2 U391 ( .A(n446), .B(n442), .Y(n182) );
  NAND2X2 U392 ( .A(n447), .B(n442), .Y(n194) );
  NAND2X2 U393 ( .A(n445), .B(n444), .Y(n176) );
  NAND2X2 U394 ( .A(n446), .B(n444), .Y(n188) );
  NAND2X2 U395 ( .A(n447), .B(n444), .Y(n200) );
  NAND2X2 U396 ( .A(n445), .B(n443), .Y(n173) );
  NAND2X2 U397 ( .A(n446), .B(n443), .Y(n185) );
  NAND2X2 U398 ( .A(n447), .B(n443), .Y(n197) );
  NAND2X2 U399 ( .A(n442), .B(n440), .Y(n158) );
  NAND2X2 U400 ( .A(n443), .B(n440), .Y(n161) );
  NAND2X2 U401 ( .A(n444), .B(n440), .Y(n164) );
  NAND2X2 U402 ( .A(n445), .B(n441), .Y(n167) );
  NAND2X2 U403 ( .A(n446), .B(n441), .Y(n179) );
  NAND2X2 U404 ( .A(n447), .B(n441), .Y(n191) );
  BUFX4 U405 ( .A(N31), .Y(n854) );
  MXI2X1 U406 ( .A(n728), .B(n729), .S0(n855), .Y(N40) );
  MX4X1 U407 ( .A(n801), .B(n799), .C(n800), .D(n798), .S0(n854), .S1(n853), 
        .Y(n728) );
  MX4X1 U408 ( .A(n797), .B(n795), .C(n796), .D(n794), .S0(n854), .S1(n853), 
        .Y(n729) );
  MXI4X1 U409 ( .A(n727), .B(n725), .C(n726), .D(n724), .S0(n852), .S1(n847), 
        .Y(n801) );
  MXI2X1 U410 ( .A(n694), .B(n695), .S0(n855), .Y(N39) );
  MX4X1 U411 ( .A(n793), .B(n791), .C(n792), .D(n790), .S0(n854), .S1(n853), 
        .Y(n694) );
  MX4X1 U412 ( .A(n789), .B(n787), .C(n788), .D(n786), .S0(n854), .S1(n853), 
        .Y(n695) );
  MXI4X1 U413 ( .A(n693), .B(n691), .C(n692), .D(n690), .S0(n852), .S1(n847), 
        .Y(n793) );
  MXI2X1 U414 ( .A(n660), .B(n661), .S0(n855), .Y(N38) );
  MX4X1 U415 ( .A(n785), .B(n783), .C(n784), .D(n782), .S0(n854), .S1(n853), 
        .Y(n660) );
  MX4X1 U416 ( .A(n781), .B(n779), .C(n780), .D(n778), .S0(n854), .S1(n853), 
        .Y(n661) );
  MXI4X1 U417 ( .A(n659), .B(n657), .C(n658), .D(n656), .S0(n851), .S1(n847), 
        .Y(n785) );
  MXI2X1 U418 ( .A(n626), .B(n627), .S0(n855), .Y(N37) );
  MX4X1 U419 ( .A(n777), .B(n775), .C(n776), .D(n774), .S0(n854), .S1(n853), 
        .Y(n626) );
  MX4X1 U420 ( .A(n773), .B(n771), .C(n772), .D(n770), .S0(n854), .S1(n853), 
        .Y(n627) );
  MXI4X1 U421 ( .A(n625), .B(n623), .C(n624), .D(n622), .S0(n850), .S1(n846), 
        .Y(n777) );
  MXI2X1 U422 ( .A(n592), .B(n593), .S0(n855), .Y(N36) );
  MX4X1 U423 ( .A(n769), .B(n767), .C(n768), .D(n766), .S0(n854), .S1(n853), 
        .Y(n592) );
  MX4X1 U424 ( .A(n765), .B(n763), .C(n764), .D(n762), .S0(n854), .S1(n853), 
        .Y(n593) );
  MXI4X1 U425 ( .A(n591), .B(n589), .C(n590), .D(n588), .S0(n850), .S1(n846), 
        .Y(n769) );
  MXI2X1 U426 ( .A(n139), .B(n140), .S0(n855), .Y(N35) );
  MX4X1 U427 ( .A(n761), .B(n759), .C(n760), .D(n758), .S0(n854), .S1(n853), 
        .Y(n139) );
  MX4X1 U428 ( .A(n757), .B(n755), .C(n756), .D(n754), .S0(n854), .S1(n853), 
        .Y(n140) );
  MXI4X1 U429 ( .A(n138), .B(n136), .C(n137), .D(n135), .S0(n850), .S1(n845), 
        .Y(n761) );
  MXI2X1 U430 ( .A(n105), .B(n106), .S0(n855), .Y(N34) );
  MX4X1 U431 ( .A(n753), .B(n751), .C(n752), .D(n750), .S0(n854), .S1(n853), 
        .Y(n105) );
  MX4X1 U432 ( .A(n749), .B(n747), .C(n748), .D(n746), .S0(n854), .S1(n853), 
        .Y(n106) );
  MXI4X1 U433 ( .A(n104), .B(n102), .C(n103), .D(n101), .S0(n848), .S1(n845), 
        .Y(n753) );
  MXI2X1 U434 ( .A(n71), .B(n72), .S0(n855), .Y(N33) );
  MX4X1 U435 ( .A(n745), .B(n743), .C(n744), .D(n742), .S0(n854), .S1(n853), 
        .Y(n71) );
  MX4X1 U436 ( .A(n741), .B(n739), .C(n740), .D(n738), .S0(n854), .S1(n853), 
        .Y(n72) );
  MXI4X1 U437 ( .A(n70), .B(n68), .C(n69), .D(n67), .S0(n848), .S1(n847), .Y(
        n745) );
  MXI2X1 U438 ( .A(n37), .B(n38), .S0(n855), .Y(N41) );
  MX4X1 U439 ( .A(n737), .B(n735), .C(n736), .D(n734), .S0(n854), .S1(n853), 
        .Y(n37) );
  MX4X1 U440 ( .A(n733), .B(n731), .C(n732), .D(n730), .S0(n854), .S1(n853), 
        .Y(n38) );
  MXI4X1 U441 ( .A(n36), .B(n34), .C(n35), .D(n33), .S0(n849), .S1(n844), .Y(
        n737) );
  BUFX4 U442 ( .A(N30), .Y(n853) );
  CLKINVX1 U443 ( .A(write_counter_count[5]), .Y(n1062) );
  CLKINVX1 U444 ( .A(write_counter_count[4]), .Y(n1061) );
  CLKINVX1 U445 ( .A(write_counter_count[0]), .Y(n985) );
  CLKBUFX3 U446 ( .A(n335), .Y(n860) );
  NAND3BX1 U447 ( .AN(write_counter_count[6]), .B(n1061), .C(
        write_counter_count[5]), .Y(n335) );
  CLKBUFX3 U448 ( .A(n154), .Y(n870) );
  NAND3X1 U449 ( .A(write_counter_count[5]), .B(write_counter_count[4]), .C(
        write_counter_count[6]), .Y(n154) );
  CLKINVX1 U450 ( .A(write_counter_count[2]), .Y(n1059) );
  CLKINVX1 U451 ( .A(write_counter_count[3]), .Y(n1060) );
  CLKINVX1 U452 ( .A(write_counter_count[1]), .Y(n1058) );
  CLKBUFX3 U453 ( .A(n302), .Y(n862) );
  NAND3BX1 U454 ( .AN(write_counter_count[6]), .B(write_counter_count[4]), .C(
        write_counter_count[5]), .Y(n302) );
  CLKBUFX3 U455 ( .A(n203), .Y(n868) );
  NAND3X1 U456 ( .A(write_counter_count[5]), .B(n1061), .C(
        write_counter_count[6]), .Y(n203) );
  CLKBUFX3 U457 ( .A(n236), .Y(n866) );
  NAND3X1 U458 ( .A(write_counter_count[4]), .B(n1062), .C(
        write_counter_count[6]), .Y(n236) );
  CLKBUFX3 U459 ( .A(n368), .Y(n858) );
  NAND3BX1 U460 ( .AN(write_counter_count[6]), .B(n1062), .C(
        write_counter_count[4]), .Y(n368) );
  CLKBUFX3 U461 ( .A(n269), .Y(n864) );
  NAND3X1 U462 ( .A(n1061), .B(n1062), .C(write_counter_count[6]), .Y(n269) );
  CLKBUFX3 U463 ( .A(n401), .Y(n856) );
  NAND3BX1 U464 ( .AN(write_counter_count[6]), .B(n1062), .C(n1061), .Y(n401)
         );
  MX4X1 U465 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .C(\mem[6][0] ), .D(
        \mem[7][0] ), .S0(n802), .S1(n843), .Y(n726) );
  MX4X1 U466 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .C(\mem[6][1] ), .D(
        \mem[7][1] ), .S0(n824), .S1(n836), .Y(n692) );
  MX4X1 U467 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .C(\mem[6][2] ), .D(
        \mem[7][2] ), .S0(n822), .S1(n841), .Y(n658) );
  MX4X1 U468 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .C(\mem[6][3] ), .D(
        \mem[7][3] ), .S0(n820), .S1(n839), .Y(n624) );
  MX4X1 U469 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .C(\mem[6][4] ), .D(
        \mem[7][4] ), .S0(n818), .S1(n838), .Y(n590) );
  MX4X1 U470 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .C(\mem[6][5] ), .D(
        \mem[7][5] ), .S0(n815), .S1(n843), .Y(n137) );
  MX4X1 U471 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .C(\mem[6][6] ), .D(
        \mem[7][6] ), .S0(n813), .S1(n836), .Y(n103) );
  MX4X1 U472 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .C(\mem[6][7] ), .D(
        \mem[7][7] ), .S0(n810), .S1(n834), .Y(n69) );
  MX4X1 U473 ( .A(valid_mem[4]), .B(valid_mem[5]), .C(valid_mem[6]), .D(
        valid_mem[7]), .S0(n808), .S1(n832), .Y(n35) );
  MX4X1 U474 ( .A(\mem[80][0] ), .B(\mem[81][0] ), .C(\mem[82][0] ), .D(
        \mem[83][0] ), .S0(n825), .S1(n827), .Y(n707) );
  MX4X1 U475 ( .A(\mem[112][0] ), .B(\mem[113][0] ), .C(\mem[114][0] ), .D(
        \mem[115][0] ), .S0(n824), .S1(n828), .Y(n699) );
  MX4X1 U476 ( .A(\mem[96][0] ), .B(\mem[97][0] ), .C(\mem[98][0] ), .D(
        \mem[99][0] ), .S0(n825), .S1(n830), .Y(n703) );
  MX4X1 U477 ( .A(\mem[64][0] ), .B(\mem[65][0] ), .C(\mem[66][0] ), .D(
        \mem[67][0] ), .S0(n825), .S1(n826), .Y(n711) );
  MX4X1 U478 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .C(\mem[18][0] ), .D(
        \mem[19][0] ), .S0(n802), .S1(n843), .Y(n723) );
  MX4X1 U479 ( .A(\mem[32][0] ), .B(\mem[33][0] ), .C(\mem[34][0] ), .D(
        \mem[35][0] ), .S0(n802), .S1(n843), .Y(n719) );
  MX4X1 U480 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .C(\mem[2][0] ), .D(
        \mem[3][0] ), .S0(n802), .S1(n843), .Y(n727) );
  MX4X1 U481 ( .A(\mem[80][1] ), .B(\mem[81][1] ), .C(\mem[82][1] ), .D(
        \mem[83][1] ), .S0(n823), .S1(n842), .Y(n673) );
  MX4X1 U482 ( .A(\mem[112][1] ), .B(\mem[113][1] ), .C(\mem[114][1] ), .D(
        \mem[115][1] ), .S0(n823), .S1(n842), .Y(n665) );
  MX4X1 U483 ( .A(\mem[96][1] ), .B(\mem[97][1] ), .C(\mem[98][1] ), .D(
        \mem[99][1] ), .S0(n823), .S1(n842), .Y(n669) );
  MX4X1 U484 ( .A(\mem[64][1] ), .B(\mem[65][1] ), .C(\mem[66][1] ), .D(
        \mem[67][1] ), .S0(n804), .S1(n826), .Y(n677) );
  MX4X1 U485 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .C(\mem[18][1] ), .D(
        \mem[19][1] ), .S0(n824), .S1(n828), .Y(n689) );
  MX4X1 U486 ( .A(\mem[48][1] ), .B(\mem[49][1] ), .C(\mem[50][1] ), .D(
        \mem[51][1] ), .S0(n803), .S1(n826), .Y(n681) );
  MX4X1 U487 ( .A(\mem[32][1] ), .B(\mem[33][1] ), .C(\mem[34][1] ), .D(
        \mem[35][1] ), .S0(n803), .S1(n829), .Y(n685) );
  MX4X1 U488 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .C(\mem[2][1] ), .D(
        \mem[3][1] ), .S0(n824), .S1(n832), .Y(n693) );
  MX4X1 U489 ( .A(\mem[80][2] ), .B(\mem[81][2] ), .C(\mem[82][2] ), .D(
        \mem[83][2] ), .S0(n821), .S1(n840), .Y(n639) );
  MX4X1 U490 ( .A(\mem[112][2] ), .B(\mem[113][2] ), .C(\mem[114][2] ), .D(
        \mem[115][2] ), .S0(n820), .S1(n839), .Y(n631) );
  MX4X1 U491 ( .A(\mem[96][2] ), .B(\mem[97][2] ), .C(\mem[98][2] ), .D(
        \mem[99][2] ), .S0(n821), .S1(n840), .Y(n635) );
  MX4X1 U492 ( .A(\mem[64][2] ), .B(\mem[65][2] ), .C(\mem[66][2] ), .D(
        \mem[67][2] ), .S0(n821), .S1(n840), .Y(n643) );
  MX4X1 U493 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .C(\mem[18][2] ), .D(
        \mem[19][2] ), .S0(n822), .S1(n841), .Y(n655) );
  MX4X1 U494 ( .A(\mem[48][2] ), .B(\mem[49][2] ), .C(\mem[50][2] ), .D(
        \mem[51][2] ), .S0(n822), .S1(n841), .Y(n647) );
  MX4X1 U495 ( .A(\mem[32][2] ), .B(\mem[33][2] ), .C(\mem[34][2] ), .D(
        \mem[35][2] ), .S0(n822), .S1(n841), .Y(n651) );
  MX4X1 U496 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .C(\mem[2][2] ), .D(
        \mem[3][2] ), .S0(n823), .S1(n842), .Y(n659) );
  MX4X1 U497 ( .A(\mem[80][3] ), .B(\mem[81][3] ), .C(\mem[82][3] ), .D(
        \mem[83][3] ), .S0(n819), .S1(n829), .Y(n605) );
  MX4X1 U498 ( .A(\mem[112][3] ), .B(\mem[113][3] ), .C(\mem[114][3] ), .D(
        \mem[115][3] ), .S0(n818), .S1(n838), .Y(n597) );
  MX4X1 U499 ( .A(\mem[96][3] ), .B(\mem[97][3] ), .C(\mem[98][3] ), .D(
        \mem[99][3] ), .S0(n818), .S1(n838), .Y(n601) );
  MX4X1 U500 ( .A(\mem[64][3] ), .B(\mem[65][3] ), .C(\mem[66][3] ), .D(
        \mem[67][3] ), .S0(n819), .S1(n827), .Y(n609) );
  MX4X1 U501 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .C(\mem[18][3] ), .D(
        \mem[19][3] ), .S0(n820), .S1(n839), .Y(n621) );
  MX4X1 U502 ( .A(\mem[48][3] ), .B(\mem[49][3] ), .C(\mem[50][3] ), .D(
        \mem[51][3] ), .S0(n819), .S1(n843), .Y(n613) );
  MX4X1 U503 ( .A(\mem[32][3] ), .B(\mem[33][3] ), .C(\mem[34][3] ), .D(
        \mem[35][3] ), .S0(n819), .S1(n828), .Y(n617) );
  MX4X1 U504 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .C(\mem[2][3] ), .D(
        \mem[3][3] ), .S0(n820), .S1(n839), .Y(n625) );
  MX4X1 U505 ( .A(\mem[80][4] ), .B(\mem[81][4] ), .C(\mem[82][4] ), .D(
        \mem[83][4] ), .S0(n816), .S1(n841), .Y(n435) );
  MX4X1 U506 ( .A(\mem[112][4] ), .B(\mem[113][4] ), .C(\mem[114][4] ), .D(
        \mem[115][4] ), .S0(n815), .S1(n828), .Y(n144) );
  MX4X1 U507 ( .A(\mem[96][4] ), .B(\mem[97][4] ), .C(\mem[98][4] ), .D(
        \mem[99][4] ), .S0(n816), .S1(n839), .Y(n148) );
  MX4X1 U508 ( .A(\mem[64][4] ), .B(\mem[65][4] ), .C(\mem[66][4] ), .D(
        \mem[67][4] ), .S0(n816), .S1(n830), .Y(n439) );
  MX4X1 U509 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .C(\mem[18][4] ), .D(
        \mem[19][4] ), .S0(n817), .S1(n837), .Y(n587) );
  MX4X1 U510 ( .A(\mem[48][4] ), .B(\mem[49][4] ), .C(\mem[50][4] ), .D(
        \mem[51][4] ), .S0(n817), .S1(n837), .Y(n579) );
  MX4X1 U511 ( .A(\mem[32][4] ), .B(\mem[33][4] ), .C(\mem[34][4] ), .D(
        \mem[35][4] ), .S0(n817), .S1(n837), .Y(n583) );
  MX4X1 U512 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .C(\mem[2][4] ), .D(
        \mem[3][4] ), .S0(n818), .S1(n838), .Y(n591) );
  MX4X1 U513 ( .A(\mem[80][5] ), .B(\mem[81][5] ), .C(\mem[82][5] ), .D(
        \mem[83][5] ), .S0(n814), .S1(n842), .Y(n118) );
  MX4X1 U514 ( .A(\mem[112][5] ), .B(\mem[113][5] ), .C(\mem[114][5] ), .D(
        \mem[115][5] ), .S0(n813), .S1(n836), .Y(n110) );
  MX4X1 U515 ( .A(\mem[96][5] ), .B(\mem[97][5] ), .C(\mem[98][5] ), .D(
        \mem[99][5] ), .S0(n813), .S1(n836), .Y(n114) );
  MX4X1 U516 ( .A(\mem[64][5] ), .B(\mem[65][5] ), .C(\mem[66][5] ), .D(
        \mem[67][5] ), .S0(n814), .S1(n826), .Y(n122) );
  MX4X1 U517 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .C(\mem[18][5] ), .D(
        \mem[19][5] ), .S0(n815), .S1(n841), .Y(n134) );
  MX4X1 U518 ( .A(\mem[48][5] ), .B(\mem[49][5] ), .C(\mem[50][5] ), .D(
        \mem[51][5] ), .S0(n814), .S1(n831), .Y(n126) );
  MX4X1 U519 ( .A(\mem[32][5] ), .B(\mem[33][5] ), .C(\mem[34][5] ), .D(
        \mem[35][5] ), .S0(n815), .S1(n842), .Y(n130) );
  MX4X1 U520 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .C(\mem[2][5] ), .D(
        \mem[3][5] ), .S0(n815), .S1(n827), .Y(n138) );
  MX4X1 U521 ( .A(\mem[80][6] ), .B(\mem[81][6] ), .C(\mem[82][6] ), .D(
        \mem[83][6] ), .S0(n811), .S1(n836), .Y(n84) );
  MX4X1 U522 ( .A(\mem[112][6] ), .B(\mem[113][6] ), .C(\mem[114][6] ), .D(
        \mem[115][6] ), .S0(n811), .S1(n837), .Y(n76) );
  MX4X1 U523 ( .A(\mem[96][6] ), .B(\mem[97][6] ), .C(\mem[98][6] ), .D(
        \mem[99][6] ), .S0(n811), .S1(n827), .Y(n80) );
  MX4X1 U524 ( .A(\mem[64][6] ), .B(\mem[65][6] ), .C(\mem[66][6] ), .D(
        \mem[67][6] ), .S0(n811), .S1(n831), .Y(n88) );
  MX4X1 U525 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .C(\mem[18][6] ), .D(
        \mem[19][6] ), .S0(n812), .S1(n835), .Y(n100) );
  MX4X1 U526 ( .A(\mem[48][6] ), .B(\mem[49][6] ), .C(\mem[50][6] ), .D(
        \mem[51][6] ), .S0(n812), .S1(n835), .Y(n92) );
  MX4X1 U527 ( .A(\mem[32][6] ), .B(\mem[33][6] ), .C(\mem[34][6] ), .D(
        \mem[35][6] ), .S0(n812), .S1(n835), .Y(n96) );
  MX4X1 U528 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .C(\mem[2][6] ), .D(
        \mem[3][6] ), .S0(n813), .S1(n836), .Y(n104) );
  MX4X1 U529 ( .A(\mem[80][7] ), .B(\mem[81][7] ), .C(\mem[82][7] ), .D(
        \mem[83][7] ), .S0(n809), .S1(n833), .Y(n50) );
  MX4X1 U530 ( .A(\mem[112][7] ), .B(\mem[113][7] ), .C(\mem[114][7] ), .D(
        \mem[115][7] ), .S0(n808), .S1(n832), .Y(n42) );
  MX4X1 U531 ( .A(\mem[96][7] ), .B(\mem[97][7] ), .C(\mem[98][7] ), .D(
        \mem[99][7] ), .S0(n808), .S1(n832), .Y(n46) );
  MX4X1 U532 ( .A(\mem[64][7] ), .B(\mem[65][7] ), .C(\mem[66][7] ), .D(
        \mem[67][7] ), .S0(n809), .S1(n833), .Y(n54) );
  MX4X1 U533 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .C(\mem[18][7] ), .D(
        \mem[19][7] ), .S0(n810), .S1(n834), .Y(n66) );
  MX4X1 U534 ( .A(\mem[48][7] ), .B(\mem[49][7] ), .C(\mem[50][7] ), .D(
        \mem[51][7] ), .S0(n809), .S1(n833), .Y(n58) );
  MX4X1 U535 ( .A(\mem[32][7] ), .B(\mem[33][7] ), .C(\mem[34][7] ), .D(
        \mem[35][7] ), .S0(n810), .S1(n834), .Y(n62) );
  MX4X1 U536 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .C(\mem[2][7] ), .D(
        \mem[3][7] ), .S0(n810), .S1(n834), .Y(n70) );
  MX4X1 U537 ( .A(valid_mem[80]), .B(valid_mem[81]), .C(valid_mem[82]), .D(
        valid_mem[83]), .S0(n806), .S1(n841), .Y(n16) );
  MX4X1 U538 ( .A(valid_mem[112]), .B(valid_mem[113]), .C(valid_mem[114]), .D(
        valid_mem[115]), .S0(n806), .S1(n832), .Y(n8) );
  MX4X1 U539 ( .A(valid_mem[96]), .B(valid_mem[97]), .C(valid_mem[98]), .D(
        valid_mem[99]), .S0(n806), .S1(n826), .Y(n12) );
  MX4X1 U540 ( .A(valid_mem[64]), .B(valid_mem[65]), .C(valid_mem[66]), .D(
        valid_mem[67]), .S0(n807), .S1(n831), .Y(n20) );
  MX4X1 U541 ( .A(valid_mem[16]), .B(valid_mem[17]), .C(valid_mem[18]), .D(
        valid_mem[19]), .S0(n807), .S1(n831), .Y(n32) );
  MX4X1 U542 ( .A(valid_mem[48]), .B(valid_mem[49]), .C(valid_mem[50]), .D(
        valid_mem[51]), .S0(n807), .S1(n831), .Y(n24) );
  MX4X1 U543 ( .A(valid_mem[32]), .B(valid_mem[33]), .C(valid_mem[34]), .D(
        valid_mem[35]), .S0(n807), .S1(n831), .Y(n28) );
  MX4X1 U544 ( .A(valid_mem[0]), .B(valid_mem[1]), .C(valid_mem[2]), .D(
        valid_mem[3]), .S0(n808), .S1(n832), .Y(n36) );
  MX4X1 U545 ( .A(\mem[56][0] ), .B(\mem[57][0] ), .C(\mem[58][0] ), .D(
        \mem[59][0] ), .S0(n825), .S1(n826), .Y(n713) );
  MX4X1 U546 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .C(\mem[10][0] ), .D(
        \mem[11][0] ), .S0(n802), .S1(n843), .Y(n725) );
  MX4X1 U547 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .C(\mem[10][1] ), .D(
        \mem[11][1] ), .S0(n824), .S1(n830), .Y(n691) );
  MX4X1 U548 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .C(\mem[10][2] ), .D(
        \mem[11][2] ), .S0(n822), .S1(n841), .Y(n657) );
  MX4X1 U549 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .C(\mem[10][3] ), .D(
        \mem[11][3] ), .S0(n820), .S1(n839), .Y(n623) );
  MX4X1 U550 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .C(\mem[10][4] ), .D(
        \mem[11][4] ), .S0(n817), .S1(n837), .Y(n589) );
  MX4X1 U551 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .C(\mem[10][5] ), .D(
        \mem[11][5] ), .S0(n815), .S1(n834), .Y(n136) );
  MX4X1 U552 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .C(\mem[10][6] ), .D(
        \mem[11][6] ), .S0(n813), .S1(n836), .Y(n102) );
  MX4X1 U553 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .C(\mem[10][7] ), .D(
        \mem[11][7] ), .S0(n810), .S1(n834), .Y(n68) );
  MX4X1 U554 ( .A(valid_mem[8]), .B(valid_mem[9]), .C(valid_mem[10]), .D(
        valid_mem[11]), .S0(n808), .S1(n832), .Y(n34) );
  MX4X1 U555 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .C(\mem[14][0] ), .D(
        \mem[15][0] ), .S0(n802), .S1(n843), .Y(n724) );
  MX4X1 U556 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .C(\mem[14][1] ), .D(
        \mem[15][1] ), .S0(n824), .S1(n835), .Y(n690) );
  MX4X1 U557 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .C(\mem[14][2] ), .D(
        \mem[15][2] ), .S0(n822), .S1(n841), .Y(n656) );
  MX4X1 U558 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .C(\mem[14][3] ), .D(
        \mem[15][3] ), .S0(n820), .S1(n839), .Y(n622) );
  MX4X1 U559 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .C(\mem[14][4] ), .D(
        \mem[15][4] ), .S0(n817), .S1(n837), .Y(n588) );
  MX4X1 U560 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .C(\mem[14][5] ), .D(
        \mem[15][5] ), .S0(n815), .S1(n840), .Y(n135) );
  MX4X1 U561 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .C(\mem[14][6] ), .D(
        \mem[15][6] ), .S0(n812), .S1(n835), .Y(n101) );
  MX4X1 U562 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .C(\mem[14][7] ), .D(
        \mem[15][7] ), .S0(n810), .S1(n834), .Y(n67) );
  MX4X1 U563 ( .A(valid_mem[12]), .B(valid_mem[13]), .C(valid_mem[14]), .D(
        valid_mem[15]), .S0(n808), .S1(n832), .Y(n33) );
  CLKBUFX3 U564 ( .A(N32), .Y(n855) );
  MXI4X1 U565 ( .A(n707), .B(n705), .C(n706), .D(n704), .S0(n852), .S1(n847), 
        .Y(n796) );
  MX4X1 U566 ( .A(\mem[92][0] ), .B(\mem[93][0] ), .C(\mem[94][0] ), .D(
        \mem[95][0] ), .S0(n825), .S1(n827), .Y(n704) );
  MX4X1 U567 ( .A(\mem[84][0] ), .B(\mem[85][0] ), .C(\mem[86][0] ), .D(
        \mem[87][0] ), .S0(n825), .S1(n826), .Y(n706) );
  MX4X1 U568 ( .A(\mem[88][0] ), .B(\mem[89][0] ), .C(\mem[90][0] ), .D(
        \mem[91][0] ), .S0(n825), .S1(n830), .Y(n705) );
  MXI4X1 U569 ( .A(n723), .B(n721), .C(n722), .D(n720), .S0(n852), .S1(n847), 
        .Y(n800) );
  MX4X1 U570 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .C(\mem[30][0] ), .D(
        \mem[31][0] ), .S0(n804), .S1(n843), .Y(n720) );
  MX4X1 U571 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .C(\mem[22][0] ), .D(
        \mem[23][0] ), .S0(n803), .S1(n843), .Y(n722) );
  MX4X1 U572 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .C(\mem[26][0] ), .D(
        \mem[27][0] ), .S0(n804), .S1(n843), .Y(n721) );
  MXI4X1 U573 ( .A(n673), .B(n671), .C(n672), .D(n670), .S0(n851), .S1(n847), 
        .Y(n788) );
  MX4X1 U574 ( .A(\mem[92][1] ), .B(\mem[93][1] ), .C(\mem[94][1] ), .D(
        \mem[95][1] ), .S0(n823), .S1(n842), .Y(n670) );
  MX4X1 U575 ( .A(\mem[84][1] ), .B(\mem[85][1] ), .C(\mem[86][1] ), .D(
        \mem[87][1] ), .S0(n823), .S1(n842), .Y(n672) );
  MX4X1 U576 ( .A(\mem[88][1] ), .B(\mem[89][1] ), .C(\mem[90][1] ), .D(
        \mem[91][1] ), .S0(n823), .S1(n842), .Y(n671) );
  MXI4X1 U577 ( .A(n689), .B(n687), .C(n688), .D(n686), .S0(n852), .S1(n847), 
        .Y(n792) );
  MX4X1 U578 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .C(\mem[30][1] ), .D(
        \mem[31][1] ), .S0(n803), .S1(n829), .Y(n686) );
  MX4X1 U579 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .C(\mem[22][1] ), .D(
        \mem[23][1] ), .S0(n824), .S1(n826), .Y(n688) );
  MX4X1 U580 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .C(\mem[26][1] ), .D(
        \mem[27][1] ), .S0(n824), .S1(n834), .Y(n687) );
  MXI4X1 U581 ( .A(n639), .B(n637), .C(n638), .D(n636), .S0(n851), .S1(n844), 
        .Y(n780) );
  MX4X1 U582 ( .A(\mem[92][2] ), .B(\mem[93][2] ), .C(\mem[94][2] ), .D(
        \mem[95][2] ), .S0(n821), .S1(n840), .Y(n636) );
  MX4X1 U583 ( .A(\mem[84][2] ), .B(\mem[85][2] ), .C(\mem[86][2] ), .D(
        \mem[87][2] ), .S0(n821), .S1(n840), .Y(n638) );
  MX4X1 U584 ( .A(\mem[88][2] ), .B(\mem[89][2] ), .C(\mem[90][2] ), .D(
        \mem[91][2] ), .S0(n821), .S1(n840), .Y(n637) );
  MXI4X1 U585 ( .A(n655), .B(n653), .C(n654), .D(n652), .S0(n851), .S1(n847), 
        .Y(n784) );
  MX4X1 U586 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .C(\mem[30][2] ), .D(
        \mem[31][2] ), .S0(n822), .S1(n841), .Y(n652) );
  MX4X1 U587 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .C(\mem[22][2] ), .D(
        \mem[23][2] ), .S0(n822), .S1(n841), .Y(n654) );
  MX4X1 U588 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .C(\mem[26][2] ), .D(
        \mem[27][2] ), .S0(n822), .S1(n841), .Y(n653) );
  MXI4X1 U589 ( .A(n605), .B(n603), .C(n604), .D(n602), .S0(n850), .S1(n846), 
        .Y(n772) );
  MX4X1 U590 ( .A(\mem[92][3] ), .B(\mem[93][3] ), .C(\mem[94][3] ), .D(
        \mem[95][3] ), .S0(n818), .S1(n838), .Y(n602) );
  MX4X1 U591 ( .A(\mem[84][3] ), .B(\mem[85][3] ), .C(\mem[86][3] ), .D(
        \mem[87][3] ), .S0(n818), .S1(n838), .Y(n604) );
  MX4X1 U592 ( .A(\mem[88][3] ), .B(\mem[89][3] ), .C(\mem[90][3] ), .D(
        \mem[91][3] ), .S0(n818), .S1(n838), .Y(n603) );
  MXI4X1 U593 ( .A(n621), .B(n619), .C(n620), .D(n618), .S0(n850), .S1(n846), 
        .Y(n776) );
  MX4X1 U594 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .C(\mem[30][3] ), .D(
        \mem[31][3] ), .S0(n820), .S1(n839), .Y(n618) );
  MX4X1 U595 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .C(\mem[22][3] ), .D(
        \mem[23][3] ), .S0(n820), .S1(n839), .Y(n620) );
  MX4X1 U596 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .C(\mem[26][3] ), .D(
        \mem[27][3] ), .S0(n820), .S1(n839), .Y(n619) );
  MXI4X1 U597 ( .A(n435), .B(n150), .C(n151), .D(n149), .S0(n851), .S1(n845), 
        .Y(n764) );
  MX4X1 U598 ( .A(\mem[92][4] ), .B(\mem[93][4] ), .C(\mem[94][4] ), .D(
        \mem[95][4] ), .S0(n816), .S1(n827), .Y(n149) );
  MX4X1 U599 ( .A(\mem[84][4] ), .B(\mem[85][4] ), .C(\mem[86][4] ), .D(
        \mem[87][4] ), .S0(n816), .S1(n831), .Y(n151) );
  MX4X1 U600 ( .A(\mem[88][4] ), .B(\mem[89][4] ), .C(\mem[90][4] ), .D(
        \mem[91][4] ), .S0(n816), .S1(n830), .Y(n150) );
  MXI4X1 U601 ( .A(n587), .B(n585), .C(n586), .D(n584), .S0(n850), .S1(n846), 
        .Y(n768) );
  MX4X1 U602 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .C(\mem[30][4] ), .D(
        \mem[31][4] ), .S0(n817), .S1(n837), .Y(n584) );
  MX4X1 U603 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .C(\mem[22][4] ), .D(
        \mem[23][4] ), .S0(n817), .S1(n837), .Y(n586) );
  MX4X1 U604 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .C(\mem[26][4] ), .D(
        \mem[27][4] ), .S0(n817), .S1(n837), .Y(n585) );
  MXI4X1 U605 ( .A(n118), .B(n116), .C(n117), .D(n115), .S0(n848), .S1(n845), 
        .Y(n756) );
  MX4X1 U606 ( .A(\mem[92][5] ), .B(\mem[93][5] ), .C(\mem[94][5] ), .D(
        \mem[95][5] ), .S0(n813), .S1(n836), .Y(n115) );
  MX4X1 U607 ( .A(\mem[84][5] ), .B(\mem[85][5] ), .C(\mem[86][5] ), .D(
        \mem[87][5] ), .S0(n814), .S1(n827), .Y(n117) );
  MX4X1 U608 ( .A(\mem[88][5] ), .B(\mem[89][5] ), .C(\mem[90][5] ), .D(
        \mem[91][5] ), .S0(n813), .S1(n836), .Y(n116) );
  MXI4X1 U609 ( .A(n134), .B(n132), .C(n133), .D(n131), .S0(n848), .S1(n845), 
        .Y(n760) );
  MX4X1 U610 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .C(\mem[30][5] ), .D(
        \mem[31][5] ), .S0(n815), .S1(n837), .Y(n131) );
  MX4X1 U611 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .C(\mem[22][5] ), .D(
        \mem[23][5] ), .S0(n815), .S1(n838), .Y(n133) );
  MX4X1 U612 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .C(\mem[26][5] ), .D(
        \mem[27][5] ), .S0(n815), .S1(n833), .Y(n132) );
  MXI4X1 U613 ( .A(n84), .B(n82), .C(n83), .D(n81), .S0(n850), .S1(n844), .Y(
        n748) );
  MX4X1 U614 ( .A(\mem[92][6] ), .B(\mem[93][6] ), .C(\mem[94][6] ), .D(
        \mem[95][6] ), .S0(n811), .S1(n829), .Y(n81) );
  MX4X1 U615 ( .A(\mem[84][6] ), .B(\mem[85][6] ), .C(\mem[86][6] ), .D(
        \mem[87][6] ), .S0(n811), .S1(n842), .Y(n83) );
  MX4X1 U616 ( .A(\mem[88][6] ), .B(\mem[89][6] ), .C(\mem[90][6] ), .D(
        \mem[91][6] ), .S0(n811), .S1(n835), .Y(n82) );
  MXI4X1 U617 ( .A(n100), .B(n98), .C(n99), .D(n97), .S0(n851), .S1(n844), .Y(
        n752) );
  MX4X1 U618 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .C(\mem[30][6] ), .D(
        \mem[31][6] ), .S0(n812), .S1(n835), .Y(n97) );
  MX4X1 U619 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .C(\mem[22][6] ), .D(
        \mem[23][6] ), .S0(n812), .S1(n835), .Y(n99) );
  MX4X1 U620 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .C(\mem[26][6] ), .D(
        \mem[27][6] ), .S0(n812), .S1(n835), .Y(n98) );
  MXI4X1 U621 ( .A(n50), .B(n48), .C(n49), .D(n47), .S0(n849), .S1(n844), .Y(
        n740) );
  MX4X1 U622 ( .A(\mem[92][7] ), .B(\mem[93][7] ), .C(\mem[94][7] ), .D(
        \mem[95][7] ), .S0(n808), .S1(n832), .Y(n47) );
  MX4X1 U623 ( .A(\mem[84][7] ), .B(\mem[85][7] ), .C(\mem[86][7] ), .D(
        \mem[87][7] ), .S0(n809), .S1(n833), .Y(n49) );
  MX4X1 U624 ( .A(\mem[88][7] ), .B(\mem[89][7] ), .C(\mem[90][7] ), .D(
        \mem[91][7] ), .S0(n809), .S1(n833), .Y(n48) );
  MXI4X1 U625 ( .A(n66), .B(n64), .C(n65), .D(n63), .S0(n848), .S1(n844), .Y(
        n744) );
  MX4X1 U626 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .C(\mem[30][7] ), .D(
        \mem[31][7] ), .S0(n810), .S1(n834), .Y(n63) );
  MX4X1 U627 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .C(\mem[22][7] ), .D(
        \mem[23][7] ), .S0(n810), .S1(n834), .Y(n65) );
  MX4X1 U628 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .C(\mem[26][7] ), .D(
        \mem[27][7] ), .S0(n810), .S1(n834), .Y(n64) );
  MXI4X1 U629 ( .A(n16), .B(n14), .C(n15), .D(n13), .S0(n849), .S1(n847), .Y(
        n732) );
  MX4X1 U630 ( .A(valid_mem[92]), .B(valid_mem[93]), .C(valid_mem[94]), .D(
        valid_mem[95]), .S0(n806), .S1(n831), .Y(n13) );
  MX4X1 U631 ( .A(valid_mem[84]), .B(valid_mem[85]), .C(valid_mem[86]), .D(
        valid_mem[87]), .S0(n806), .S1(n826), .Y(n15) );
  MX4X1 U632 ( .A(valid_mem[88]), .B(valid_mem[89]), .C(valid_mem[90]), .D(
        valid_mem[91]), .S0(n806), .S1(n833), .Y(n14) );
  MXI4X1 U633 ( .A(n32), .B(n30), .C(n31), .D(n29), .S0(n849), .S1(n844), .Y(
        n736) );
  MX4X1 U634 ( .A(valid_mem[28]), .B(valid_mem[29]), .C(valid_mem[30]), .D(
        valid_mem[31]), .S0(n807), .S1(n831), .Y(n29) );
  MX4X1 U635 ( .A(valid_mem[20]), .B(valid_mem[21]), .C(valid_mem[22]), .D(
        valid_mem[23]), .S0(n807), .S1(n831), .Y(n31) );
  MX4X1 U636 ( .A(valid_mem[24]), .B(valid_mem[25]), .C(valid_mem[26]), .D(
        valid_mem[27]), .S0(n807), .S1(n831), .Y(n30) );
  MXI4X1 U637 ( .A(n711), .B(n709), .C(n710), .D(n708), .S0(n852), .S1(n847), 
        .Y(n797) );
  MX4X1 U638 ( .A(\mem[76][0] ), .B(\mem[77][0] ), .C(\mem[78][0] ), .D(
        \mem[79][0] ), .S0(n825), .S1(n826), .Y(n708) );
  MX4X1 U639 ( .A(\mem[68][0] ), .B(\mem[69][0] ), .C(\mem[70][0] ), .D(
        \mem[71][0] ), .S0(n825), .S1(n828), .Y(n710) );
  MX4X1 U640 ( .A(\mem[72][0] ), .B(\mem[73][0] ), .C(\mem[74][0] ), .D(
        \mem[75][0] ), .S0(n825), .S1(n826), .Y(n709) );
  MXI4X1 U641 ( .A(n677), .B(n675), .C(n676), .D(n674), .S0(n851), .S1(n847), 
        .Y(n789) );
  MX4X1 U642 ( .A(\mem[76][1] ), .B(\mem[77][1] ), .C(\mem[78][1] ), .D(
        \mem[79][1] ), .S0(n805), .S1(n826), .Y(n674) );
  MX4X1 U643 ( .A(\mem[68][1] ), .B(\mem[69][1] ), .C(\mem[70][1] ), .D(
        \mem[71][1] ), .S0(n803), .S1(n829), .Y(n676) );
  MX4X1 U644 ( .A(\mem[72][1] ), .B(\mem[73][1] ), .C(\mem[74][1] ), .D(
        \mem[75][1] ), .S0(n804), .S1(n841), .Y(n675) );
  MXI4X1 U645 ( .A(n643), .B(n641), .C(n642), .D(n640), .S0(n851), .S1(n846), 
        .Y(n781) );
  MX4X1 U646 ( .A(\mem[76][2] ), .B(\mem[77][2] ), .C(\mem[78][2] ), .D(
        \mem[79][2] ), .S0(n821), .S1(n840), .Y(n640) );
  MX4X1 U647 ( .A(\mem[68][2] ), .B(\mem[69][2] ), .C(\mem[70][2] ), .D(
        \mem[71][2] ), .S0(n821), .S1(n840), .Y(n642) );
  MX4X1 U648 ( .A(\mem[72][2] ), .B(\mem[73][2] ), .C(\mem[74][2] ), .D(
        \mem[75][2] ), .S0(n821), .S1(n840), .Y(n641) );
  MXI4X1 U649 ( .A(n609), .B(n607), .C(n608), .D(n606), .S0(n850), .S1(n846), 
        .Y(n773) );
  MX4X1 U650 ( .A(\mem[76][3] ), .B(\mem[77][3] ), .C(\mem[78][3] ), .D(
        \mem[79][3] ), .S0(n819), .S1(n832), .Y(n606) );
  MX4X1 U651 ( .A(\mem[68][3] ), .B(\mem[69][3] ), .C(\mem[70][3] ), .D(
        \mem[71][3] ), .S0(n819), .S1(n828), .Y(n608) );
  MX4X1 U652 ( .A(\mem[72][3] ), .B(\mem[73][3] ), .C(\mem[74][3] ), .D(
        \mem[75][3] ), .S0(n819), .S1(n836), .Y(n607) );
  MXI4X1 U653 ( .A(n439), .B(n437), .C(n438), .D(n436), .S0(n848), .S1(n845), 
        .Y(n765) );
  MX4X1 U654 ( .A(\mem[76][4] ), .B(\mem[77][4] ), .C(\mem[78][4] ), .D(
        \mem[79][4] ), .S0(n816), .S1(n838), .Y(n436) );
  MX4X1 U655 ( .A(\mem[68][4] ), .B(\mem[69][4] ), .C(\mem[70][4] ), .D(
        \mem[71][4] ), .S0(n816), .S1(n828), .Y(n438) );
  MX4X1 U656 ( .A(\mem[72][4] ), .B(\mem[73][4] ), .C(\mem[74][4] ), .D(
        \mem[75][4] ), .S0(n816), .S1(n840), .Y(n437) );
  MXI4X1 U657 ( .A(n122), .B(n120), .C(n121), .D(n119), .S0(n849), .S1(n845), 
        .Y(n757) );
  MX4X1 U658 ( .A(\mem[76][5] ), .B(\mem[77][5] ), .C(\mem[78][5] ), .D(
        \mem[79][5] ), .S0(n814), .S1(n828), .Y(n119) );
  MX4X1 U659 ( .A(\mem[68][5] ), .B(\mem[69][5] ), .C(\mem[70][5] ), .D(
        \mem[71][5] ), .S0(n814), .S1(n827), .Y(n121) );
  MX4X1 U660 ( .A(\mem[72][5] ), .B(\mem[73][5] ), .C(\mem[74][5] ), .D(
        \mem[75][5] ), .S0(n814), .S1(n840), .Y(n120) );
  MXI4X1 U661 ( .A(n88), .B(n86), .C(n87), .D(n85), .S0(n848), .S1(n844), .Y(
        n749) );
  MX4X1 U662 ( .A(\mem[76][6] ), .B(\mem[77][6] ), .C(\mem[78][6] ), .D(
        \mem[79][6] ), .S0(n811), .S1(n828), .Y(n85) );
  MX4X1 U663 ( .A(\mem[68][6] ), .B(\mem[69][6] ), .C(\mem[70][6] ), .D(
        \mem[71][6] ), .S0(n811), .S1(n827), .Y(n87) );
  MX4X1 U664 ( .A(\mem[72][6] ), .B(\mem[73][6] ), .C(\mem[74][6] ), .D(
        \mem[75][6] ), .S0(n811), .S1(n836), .Y(n86) );
  MXI4X1 U665 ( .A(n54), .B(n52), .C(n53), .D(n51), .S0(n849), .S1(N28), .Y(
        n741) );
  MX4X1 U666 ( .A(\mem[76][7] ), .B(\mem[77][7] ), .C(\mem[78][7] ), .D(
        \mem[79][7] ), .S0(n809), .S1(n833), .Y(n51) );
  MX4X1 U667 ( .A(\mem[68][7] ), .B(\mem[69][7] ), .C(\mem[70][7] ), .D(
        \mem[71][7] ), .S0(n809), .S1(n833), .Y(n53) );
  MX4X1 U668 ( .A(\mem[72][7] ), .B(\mem[73][7] ), .C(\mem[74][7] ), .D(
        \mem[75][7] ), .S0(n809), .S1(n833), .Y(n52) );
  MXI4X1 U669 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n849), .S1(n844), .Y(
        n733) );
  MX4X1 U670 ( .A(valid_mem[76]), .B(valid_mem[77]), .C(valid_mem[78]), .D(
        valid_mem[79]), .S0(n806), .S1(n835), .Y(n17) );
  MX4X1 U671 ( .A(valid_mem[68]), .B(valid_mem[69]), .C(valid_mem[70]), .D(
        valid_mem[71]), .S0(n806), .S1(n826), .Y(n19) );
  MX4X1 U672 ( .A(valid_mem[72]), .B(valid_mem[73]), .C(valid_mem[74]), .D(
        valid_mem[75]), .S0(n806), .S1(n837), .Y(n18) );
  MXI4X1 U673 ( .A(n699), .B(n697), .C(n698), .D(n696), .S0(n852), .S1(n847), 
        .Y(n794) );
  MX4X1 U674 ( .A(\mem[124][0] ), .B(\mem[125][0] ), .C(\mem[126][0] ), .D(
        \mem[127][0] ), .S0(n824), .S1(n827), .Y(n696) );
  MX4X1 U675 ( .A(\mem[116][0] ), .B(\mem[117][0] ), .C(\mem[118][0] ), .D(
        \mem[119][0] ), .S0(n824), .S1(n828), .Y(n698) );
  MX4X1 U676 ( .A(\mem[120][0] ), .B(\mem[121][0] ), .C(\mem[122][0] ), .D(
        \mem[123][0] ), .S0(n824), .S1(n839), .Y(n697) );
  MXI4X1 U677 ( .A(n715), .B(n713), .C(n714), .D(n712), .S0(n852), .S1(n847), 
        .Y(n798) );
  MX4X1 U678 ( .A(\mem[60][0] ), .B(\mem[61][0] ), .C(\mem[62][0] ), .D(
        \mem[63][0] ), .S0(n825), .S1(n830), .Y(n712) );
  MX4X1 U679 ( .A(\mem[52][0] ), .B(\mem[53][0] ), .C(\mem[54][0] ), .D(
        \mem[55][0] ), .S0(n825), .S1(n830), .Y(n714) );
  MX4X1 U680 ( .A(\mem[48][0] ), .B(\mem[49][0] ), .C(\mem[50][0] ), .D(
        \mem[51][0] ), .S0(n804), .S1(n843), .Y(n715) );
  MXI4X1 U681 ( .A(n665), .B(n663), .C(n664), .D(n662), .S0(n851), .S1(n846), 
        .Y(n786) );
  MX4X1 U682 ( .A(\mem[124][1] ), .B(\mem[125][1] ), .C(\mem[126][1] ), .D(
        \mem[127][1] ), .S0(n823), .S1(n842), .Y(n662) );
  MX4X1 U683 ( .A(\mem[116][1] ), .B(\mem[117][1] ), .C(\mem[118][1] ), .D(
        \mem[119][1] ), .S0(n823), .S1(n842), .Y(n664) );
  MX4X1 U684 ( .A(\mem[120][1] ), .B(\mem[121][1] ), .C(\mem[122][1] ), .D(
        \mem[123][1] ), .S0(n823), .S1(n842), .Y(n663) );
  MXI4X1 U685 ( .A(n681), .B(n679), .C(n680), .D(n678), .S0(n852), .S1(n847), 
        .Y(n790) );
  MX4X1 U686 ( .A(\mem[60][1] ), .B(\mem[61][1] ), .C(\mem[62][1] ), .D(
        \mem[63][1] ), .S0(n804), .S1(n830), .Y(n678) );
  MX4X1 U687 ( .A(\mem[52][1] ), .B(\mem[53][1] ), .C(\mem[54][1] ), .D(
        \mem[55][1] ), .S0(n802), .S1(n829), .Y(n680) );
  MX4X1 U688 ( .A(\mem[56][1] ), .B(\mem[57][1] ), .C(\mem[58][1] ), .D(
        \mem[59][1] ), .S0(n803), .S1(n827), .Y(n679) );
  MXI4X1 U689 ( .A(n631), .B(n629), .C(n630), .D(n628), .S0(n851), .S1(n845), 
        .Y(n778) );
  MX4X1 U690 ( .A(\mem[124][2] ), .B(\mem[125][2] ), .C(\mem[126][2] ), .D(
        \mem[127][2] ), .S0(n820), .S1(n839), .Y(n628) );
  MX4X1 U691 ( .A(\mem[116][2] ), .B(\mem[117][2] ), .C(\mem[118][2] ), .D(
        \mem[119][2] ), .S0(n820), .S1(n839), .Y(n630) );
  MX4X1 U692 ( .A(\mem[120][2] ), .B(\mem[121][2] ), .C(\mem[122][2] ), .D(
        \mem[123][2] ), .S0(n820), .S1(n839), .Y(n629) );
  MXI4X1 U693 ( .A(n647), .B(n645), .C(n646), .D(n644), .S0(n851), .S1(n845), 
        .Y(n782) );
  MX4X1 U694 ( .A(\mem[60][2] ), .B(\mem[61][2] ), .C(\mem[62][2] ), .D(
        \mem[63][2] ), .S0(n821), .S1(n840), .Y(n644) );
  MX4X1 U695 ( .A(\mem[52][2] ), .B(\mem[53][2] ), .C(\mem[54][2] ), .D(
        \mem[55][2] ), .S0(n822), .S1(n841), .Y(n646) );
  MX4X1 U696 ( .A(\mem[56][2] ), .B(\mem[57][2] ), .C(\mem[58][2] ), .D(
        \mem[59][2] ), .S0(n821), .S1(n840), .Y(n645) );
  MXI4X1 U697 ( .A(n597), .B(n595), .C(n596), .D(n594), .S0(n850), .S1(n846), 
        .Y(n770) );
  MX4X1 U698 ( .A(\mem[124][3] ), .B(\mem[125][3] ), .C(\mem[126][3] ), .D(
        \mem[127][3] ), .S0(n818), .S1(n838), .Y(n594) );
  MX4X1 U699 ( .A(\mem[116][3] ), .B(\mem[117][3] ), .C(\mem[118][3] ), .D(
        \mem[119][3] ), .S0(n818), .S1(n838), .Y(n596) );
  MX4X1 U700 ( .A(\mem[120][3] ), .B(\mem[121][3] ), .C(\mem[122][3] ), .D(
        \mem[123][3] ), .S0(n818), .S1(n838), .Y(n595) );
  MXI4X1 U701 ( .A(n613), .B(n611), .C(n612), .D(n610), .S0(n850), .S1(n846), 
        .Y(n774) );
  MX4X1 U702 ( .A(\mem[60][3] ), .B(\mem[61][3] ), .C(\mem[62][3] ), .D(
        \mem[63][3] ), .S0(n819), .S1(n829), .Y(n610) );
  MX4X1 U703 ( .A(\mem[52][3] ), .B(\mem[53][3] ), .C(\mem[54][3] ), .D(
        \mem[55][3] ), .S0(n819), .S1(n828), .Y(n612) );
  MX4X1 U704 ( .A(\mem[56][3] ), .B(\mem[57][3] ), .C(\mem[58][3] ), .D(
        \mem[59][3] ), .S0(n819), .S1(n829), .Y(n611) );
  MXI4X1 U705 ( .A(n144), .B(n142), .C(n143), .D(n141), .S0(n850), .S1(n845), 
        .Y(n762) );
  MX4X1 U706 ( .A(\mem[124][4] ), .B(\mem[125][4] ), .C(\mem[126][4] ), .D(
        \mem[127][4] ), .S0(n815), .S1(n828), .Y(n141) );
  MX4X1 U707 ( .A(\mem[116][4] ), .B(\mem[117][4] ), .C(\mem[118][4] ), .D(
        \mem[119][4] ), .S0(n815), .S1(n829), .Y(n143) );
  MX4X1 U708 ( .A(\mem[120][4] ), .B(\mem[121][4] ), .C(\mem[122][4] ), .D(
        \mem[123][4] ), .S0(n815), .S1(n827), .Y(n142) );
  MXI4X1 U709 ( .A(n579), .B(n577), .C(n578), .D(n576), .S0(n850), .S1(n846), 
        .Y(n766) );
  MX4X1 U710 ( .A(\mem[60][4] ), .B(\mem[61][4] ), .C(\mem[62][4] ), .D(
        \mem[63][4] ), .S0(n816), .S1(n834), .Y(n576) );
  MX4X1 U711 ( .A(\mem[52][4] ), .B(\mem[53][4] ), .C(\mem[54][4] ), .D(
        \mem[55][4] ), .S0(n817), .S1(n837), .Y(n578) );
  MX4X1 U712 ( .A(\mem[56][4] ), .B(\mem[57][4] ), .C(\mem[58][4] ), .D(
        \mem[59][4] ), .S0(n817), .S1(n837), .Y(n577) );
  MXI4X1 U713 ( .A(n110), .B(n108), .C(n109), .D(n107), .S0(n852), .S1(n845), 
        .Y(n754) );
  MX4X1 U714 ( .A(\mem[124][5] ), .B(\mem[125][5] ), .C(\mem[126][5] ), .D(
        \mem[127][5] ), .S0(n813), .S1(n836), .Y(n107) );
  MX4X1 U715 ( .A(\mem[116][5] ), .B(\mem[117][5] ), .C(\mem[118][5] ), .D(
        \mem[119][5] ), .S0(n813), .S1(n836), .Y(n109) );
  MX4X1 U716 ( .A(\mem[120][5] ), .B(\mem[121][5] ), .C(\mem[122][5] ), .D(
        \mem[123][5] ), .S0(n813), .S1(n836), .Y(n108) );
  MXI4X1 U717 ( .A(n126), .B(n124), .C(n125), .D(n123), .S0(n848), .S1(n845), 
        .Y(n758) );
  MX4X1 U718 ( .A(\mem[60][5] ), .B(\mem[61][5] ), .C(\mem[62][5] ), .D(
        \mem[63][5] ), .S0(n814), .S1(n840), .Y(n123) );
  MX4X1 U719 ( .A(\mem[52][5] ), .B(\mem[53][5] ), .C(\mem[54][5] ), .D(
        \mem[55][5] ), .S0(n814), .S1(n832), .Y(n125) );
  MX4X1 U720 ( .A(\mem[56][5] ), .B(\mem[57][5] ), .C(\mem[58][5] ), .D(
        \mem[59][5] ), .S0(n814), .S1(n839), .Y(n124) );
  MXI4X1 U721 ( .A(n76), .B(n74), .C(n75), .D(n73), .S0(n849), .S1(n844), .Y(
        n746) );
  MX4X1 U722 ( .A(\mem[124][6] ), .B(\mem[125][6] ), .C(\mem[126][6] ), .D(
        \mem[127][6] ), .S0(n810), .S1(n834), .Y(n73) );
  MX4X1 U723 ( .A(\mem[116][6] ), .B(\mem[117][6] ), .C(\mem[118][6] ), .D(
        \mem[119][6] ), .S0(n810), .S1(n834), .Y(n75) );
  MX4X1 U724 ( .A(\mem[120][6] ), .B(\mem[121][6] ), .C(\mem[122][6] ), .D(
        \mem[123][6] ), .S0(n810), .S1(n834), .Y(n74) );
  MXI4X1 U725 ( .A(n92), .B(n90), .C(n91), .D(n89), .S0(n848), .S1(n844), .Y(
        n750) );
  MX4X1 U726 ( .A(\mem[60][6] ), .B(\mem[61][6] ), .C(\mem[62][6] ), .D(
        \mem[63][6] ), .S0(n812), .S1(n835), .Y(n89) );
  MX4X1 U727 ( .A(\mem[52][6] ), .B(\mem[53][6] ), .C(\mem[54][6] ), .D(
        \mem[55][6] ), .S0(n812), .S1(n835), .Y(n91) );
  MX4X1 U728 ( .A(\mem[56][6] ), .B(\mem[57][6] ), .C(\mem[58][6] ), .D(
        \mem[59][6] ), .S0(n812), .S1(n835), .Y(n90) );
  MXI4X1 U729 ( .A(n42), .B(n40), .C(n41), .D(n39), .S0(n849), .S1(n846), .Y(
        n738) );
  MX4X1 U730 ( .A(\mem[124][7] ), .B(\mem[125][7] ), .C(\mem[126][7] ), .D(
        \mem[127][7] ), .S0(n808), .S1(n832), .Y(n39) );
  MX4X1 U731 ( .A(\mem[116][7] ), .B(\mem[117][7] ), .C(\mem[118][7] ), .D(
        \mem[119][7] ), .S0(n808), .S1(n832), .Y(n41) );
  MX4X1 U732 ( .A(\mem[120][7] ), .B(\mem[121][7] ), .C(\mem[122][7] ), .D(
        \mem[123][7] ), .S0(n808), .S1(n832), .Y(n40) );
  MXI4X1 U733 ( .A(n58), .B(n56), .C(n57), .D(n55), .S0(n852), .S1(n844), .Y(
        n742) );
  MX4X1 U734 ( .A(\mem[60][7] ), .B(\mem[61][7] ), .C(\mem[62][7] ), .D(
        \mem[63][7] ), .S0(n809), .S1(n833), .Y(n55) );
  MX4X1 U735 ( .A(\mem[52][7] ), .B(\mem[53][7] ), .C(\mem[54][7] ), .D(
        \mem[55][7] ), .S0(n809), .S1(n833), .Y(n57) );
  MX4X1 U736 ( .A(\mem[56][7] ), .B(\mem[57][7] ), .C(\mem[58][7] ), .D(
        \mem[59][7] ), .S0(n809), .S1(n833), .Y(n56) );
  MXI4X1 U737 ( .A(n8), .B(n6), .C(n7), .D(n5), .S0(n849), .S1(n845), .Y(n730)
         );
  MX4X1 U738 ( .A(valid_mem[124]), .B(valid_mem[125]), .C(valid_mem[126]), .D(
        valid_mem[127]), .S0(n802), .S1(n827), .Y(n5) );
  MX4X1 U739 ( .A(valid_mem[120]), .B(valid_mem[121]), .C(valid_mem[122]), .D(
        valid_mem[123]), .S0(n805), .S1(n843), .Y(n6) );
  MX4X1 U740 ( .A(valid_mem[116]), .B(valid_mem[117]), .C(valid_mem[118]), .D(
        valid_mem[119]), .S0(n806), .S1(n834), .Y(n7) );
  MXI4X1 U741 ( .A(n24), .B(n22), .C(n23), .D(n21), .S0(n849), .S1(n846), .Y(
        n734) );
  MX4X1 U742 ( .A(valid_mem[60]), .B(valid_mem[61]), .C(valid_mem[62]), .D(
        valid_mem[63]), .S0(n807), .S1(n831), .Y(n21) );
  MX4X1 U743 ( .A(valid_mem[52]), .B(valid_mem[53]), .C(valid_mem[54]), .D(
        valid_mem[55]), .S0(n807), .S1(n831), .Y(n23) );
  MX4X1 U744 ( .A(valid_mem[56]), .B(valid_mem[57]), .C(valid_mem[58]), .D(
        valid_mem[59]), .S0(n807), .S1(n831), .Y(n22) );
  NAND2X1 U745 ( .A(n165), .B(n166), .Y(n452) );
  OAI21XL U746 ( .A0(n870), .A1(n167), .B0(valid_mem[123]), .Y(n166) );
  NAND2X1 U747 ( .A(n168), .B(n169), .Y(n453) );
  OAI21XL U748 ( .A0(n870), .A1(n170), .B0(valid_mem[122]), .Y(n169) );
  NAND2X1 U749 ( .A(n171), .B(n172), .Y(n454) );
  OAI21XL U750 ( .A0(n870), .A1(n173), .B0(valid_mem[121]), .Y(n172) );
  NAND2X1 U751 ( .A(n174), .B(n175), .Y(n455) );
  OAI21XL U752 ( .A0(n870), .A1(n176), .B0(valid_mem[120]), .Y(n175) );
  NAND2X1 U753 ( .A(n177), .B(n178), .Y(n456) );
  OAI21XL U754 ( .A0(n870), .A1(n179), .B0(valid_mem[119]), .Y(n178) );
  NAND2X1 U755 ( .A(n180), .B(n181), .Y(n457) );
  OAI21XL U756 ( .A0(n870), .A1(n182), .B0(valid_mem[118]), .Y(n181) );
  NAND2X1 U757 ( .A(n183), .B(n184), .Y(n458) );
  OAI21XL U758 ( .A0(n870), .A1(n185), .B0(valid_mem[117]), .Y(n184) );
  NAND2X1 U759 ( .A(n186), .B(n187), .Y(n459) );
  OAI21XL U760 ( .A0(n870), .A1(n188), .B0(valid_mem[116]), .Y(n187) );
  NAND2X1 U761 ( .A(n189), .B(n190), .Y(n460) );
  OAI21XL U762 ( .A0(n870), .A1(n191), .B0(valid_mem[115]), .Y(n190) );
  NAND2X1 U763 ( .A(n192), .B(n193), .Y(n461) );
  OAI21XL U764 ( .A0(n870), .A1(n194), .B0(valid_mem[114]), .Y(n193) );
  NAND2X1 U765 ( .A(n195), .B(n196), .Y(n462) );
  OAI21XL U766 ( .A0(n870), .A1(n197), .B0(valid_mem[113]), .Y(n196) );
  NAND2X1 U767 ( .A(n198), .B(n199), .Y(n463) );
  OAI21XL U768 ( .A0(n870), .A1(n200), .B0(valid_mem[112]), .Y(n199) );
  NAND2X1 U769 ( .A(n156), .B(n157), .Y(n449) );
  OAI21XL U770 ( .A0(n870), .A1(n158), .B0(valid_mem[126]), .Y(n157) );
  NAND2X1 U771 ( .A(n159), .B(n160), .Y(n450) );
  OAI21XL U772 ( .A0(n870), .A1(n161), .B0(valid_mem[125]), .Y(n160) );
  NAND2X1 U773 ( .A(n162), .B(n163), .Y(n451) );
  OAI21XL U774 ( .A0(n870), .A1(n164), .B0(valid_mem[124]), .Y(n163) );
  MXI4X1 U775 ( .A(n703), .B(n701), .C(n702), .D(n700), .S0(n852), .S1(n847), 
        .Y(n795) );
  MX4X1 U776 ( .A(\mem[108][0] ), .B(\mem[109][0] ), .C(\mem[110][0] ), .D(
        \mem[111][0] ), .S0(n824), .S1(n833), .Y(n700) );
  MX4X1 U777 ( .A(\mem[100][0] ), .B(\mem[101][0] ), .C(\mem[102][0] ), .D(
        \mem[103][0] ), .S0(n825), .S1(n826), .Y(n702) );
  MX4X1 U778 ( .A(\mem[104][0] ), .B(\mem[105][0] ), .C(\mem[106][0] ), .D(
        \mem[107][0] ), .S0(n824), .S1(n837), .Y(n701) );
  MXI4X1 U779 ( .A(n719), .B(n717), .C(n718), .D(n716), .S0(n852), .S1(n847), 
        .Y(n799) );
  MX4X1 U780 ( .A(\mem[44][0] ), .B(\mem[45][0] ), .C(\mem[46][0] ), .D(
        \mem[47][0] ), .S0(n803), .S1(n843), .Y(n716) );
  MX4X1 U781 ( .A(\mem[36][0] ), .B(\mem[37][0] ), .C(\mem[38][0] ), .D(
        \mem[39][0] ), .S0(n802), .S1(n843), .Y(n718) );
  MX4X1 U782 ( .A(\mem[40][0] ), .B(\mem[41][0] ), .C(\mem[42][0] ), .D(
        \mem[43][0] ), .S0(n804), .S1(n843), .Y(n717) );
  MXI4X1 U783 ( .A(n669), .B(n667), .C(n668), .D(n666), .S0(n851), .S1(n846), 
        .Y(n787) );
  MX4X1 U784 ( .A(\mem[108][1] ), .B(\mem[109][1] ), .C(\mem[110][1] ), .D(
        \mem[111][1] ), .S0(n823), .S1(n842), .Y(n666) );
  MX4X1 U785 ( .A(\mem[100][1] ), .B(\mem[101][1] ), .C(\mem[102][1] ), .D(
        \mem[103][1] ), .S0(n823), .S1(n842), .Y(n668) );
  MX4X1 U786 ( .A(\mem[104][1] ), .B(\mem[105][1] ), .C(\mem[106][1] ), .D(
        \mem[107][1] ), .S0(n823), .S1(n842), .Y(n667) );
  MXI4X1 U787 ( .A(n685), .B(n683), .C(n684), .D(n682), .S0(n852), .S1(n847), 
        .Y(n791) );
  MX4X1 U788 ( .A(\mem[44][1] ), .B(\mem[45][1] ), .C(\mem[46][1] ), .D(
        \mem[47][1] ), .S0(n802), .S1(n826), .Y(n682) );
  MX4X1 U789 ( .A(\mem[36][1] ), .B(\mem[37][1] ), .C(\mem[38][1] ), .D(
        \mem[39][1] ), .S0(n802), .S1(n829), .Y(n684) );
  MX4X1 U790 ( .A(\mem[40][1] ), .B(\mem[41][1] ), .C(\mem[42][1] ), .D(
        \mem[43][1] ), .S0(n804), .S1(n829), .Y(n683) );
  MXI4X1 U791 ( .A(n635), .B(n633), .C(n634), .D(n632), .S0(n851), .S1(n845), 
        .Y(n779) );
  MX4X1 U792 ( .A(\mem[108][2] ), .B(\mem[109][2] ), .C(\mem[110][2] ), .D(
        \mem[111][2] ), .S0(n820), .S1(n839), .Y(n632) );
  MX4X1 U793 ( .A(\mem[100][2] ), .B(\mem[101][2] ), .C(\mem[102][2] ), .D(
        \mem[103][2] ), .S0(n821), .S1(n840), .Y(n634) );
  MX4X1 U794 ( .A(\mem[104][2] ), .B(\mem[105][2] ), .C(\mem[106][2] ), .D(
        \mem[107][2] ), .S0(n821), .S1(n840), .Y(n633) );
  MXI4X1 U795 ( .A(n651), .B(n649), .C(n650), .D(n648), .S0(n851), .S1(n845), 
        .Y(n783) );
  MX4X1 U796 ( .A(\mem[44][2] ), .B(\mem[45][2] ), .C(\mem[46][2] ), .D(
        \mem[47][2] ), .S0(n822), .S1(n841), .Y(n648) );
  MX4X1 U797 ( .A(\mem[36][2] ), .B(\mem[37][2] ), .C(\mem[38][2] ), .D(
        \mem[39][2] ), .S0(n822), .S1(n841), .Y(n650) );
  MX4X1 U798 ( .A(\mem[40][2] ), .B(\mem[41][2] ), .C(\mem[42][2] ), .D(
        \mem[43][2] ), .S0(n822), .S1(n841), .Y(n649) );
  MXI4X1 U799 ( .A(n601), .B(n599), .C(n600), .D(n598), .S0(n850), .S1(n846), 
        .Y(n771) );
  MX4X1 U800 ( .A(\mem[108][3] ), .B(\mem[109][3] ), .C(\mem[110][3] ), .D(
        \mem[111][3] ), .S0(n818), .S1(n838), .Y(n598) );
  MX4X1 U801 ( .A(\mem[100][3] ), .B(\mem[101][3] ), .C(\mem[102][3] ), .D(
        \mem[103][3] ), .S0(n818), .S1(n838), .Y(n600) );
  MX4X1 U802 ( .A(\mem[104][3] ), .B(\mem[105][3] ), .C(\mem[106][3] ), .D(
        \mem[107][3] ), .S0(n818), .S1(n838), .Y(n599) );
  MXI4X1 U803 ( .A(n617), .B(n615), .C(n616), .D(n614), .S0(n850), .S1(n846), 
        .Y(n775) );
  MX4X1 U804 ( .A(\mem[44][3] ), .B(\mem[45][3] ), .C(\mem[46][3] ), .D(
        \mem[47][3] ), .S0(n819), .S1(n830), .Y(n614) );
  MX4X1 U805 ( .A(\mem[36][3] ), .B(\mem[37][3] ), .C(\mem[38][3] ), .D(
        \mem[39][3] ), .S0(n819), .S1(n830), .Y(n616) );
  MX4X1 U806 ( .A(\mem[40][3] ), .B(\mem[41][3] ), .C(\mem[42][3] ), .D(
        \mem[43][3] ), .S0(n819), .S1(n827), .Y(n615) );
  MXI4X1 U807 ( .A(n148), .B(n146), .C(n147), .D(n145), .S0(n848), .S1(n845), 
        .Y(n763) );
  MX4X1 U808 ( .A(\mem[108][4] ), .B(\mem[109][4] ), .C(\mem[110][4] ), .D(
        \mem[111][4] ), .S0(n816), .S1(n829), .Y(n145) );
  MX4X1 U809 ( .A(\mem[100][4] ), .B(\mem[101][4] ), .C(\mem[102][4] ), .D(
        \mem[103][4] ), .S0(n816), .S1(n830), .Y(n147) );
  MX4X1 U810 ( .A(\mem[104][4] ), .B(\mem[105][4] ), .C(\mem[106][4] ), .D(
        \mem[107][4] ), .S0(n816), .S1(n833), .Y(n146) );
  MXI4X1 U811 ( .A(n583), .B(n581), .C(n582), .D(n580), .S0(n850), .S1(n846), 
        .Y(n767) );
  MX4X1 U812 ( .A(\mem[44][4] ), .B(\mem[45][4] ), .C(\mem[46][4] ), .D(
        \mem[47][4] ), .S0(n817), .S1(n837), .Y(n580) );
  MX4X1 U813 ( .A(\mem[36][4] ), .B(\mem[37][4] ), .C(\mem[38][4] ), .D(
        \mem[39][4] ), .S0(n817), .S1(n837), .Y(n582) );
  MX4X1 U814 ( .A(\mem[40][4] ), .B(\mem[41][4] ), .C(\mem[42][4] ), .D(
        \mem[43][4] ), .S0(n817), .S1(n837), .Y(n581) );
  MXI4X1 U815 ( .A(n114), .B(n112), .C(n113), .D(n111), .S0(n848), .S1(n845), 
        .Y(n755) );
  MX4X1 U816 ( .A(\mem[108][5] ), .B(\mem[109][5] ), .C(\mem[110][5] ), .D(
        \mem[111][5] ), .S0(n813), .S1(n836), .Y(n111) );
  MX4X1 U817 ( .A(\mem[100][5] ), .B(\mem[101][5] ), .C(\mem[102][5] ), .D(
        \mem[103][5] ), .S0(n813), .S1(n836), .Y(n113) );
  MX4X1 U818 ( .A(\mem[104][5] ), .B(\mem[105][5] ), .C(\mem[106][5] ), .D(
        \mem[107][5] ), .S0(n813), .S1(n836), .Y(n112) );
  MXI4X1 U819 ( .A(n130), .B(n128), .C(n129), .D(n127), .S0(n851), .S1(n845), 
        .Y(n759) );
  MX4X1 U820 ( .A(\mem[44][5] ), .B(\mem[45][5] ), .C(\mem[46][5] ), .D(
        \mem[47][5] ), .S0(n814), .S1(n843), .Y(n127) );
  MX4X1 U821 ( .A(\mem[36][5] ), .B(\mem[37][5] ), .C(\mem[38][5] ), .D(
        \mem[39][5] ), .S0(n814), .S1(n839), .Y(n129) );
  MX4X1 U822 ( .A(\mem[40][5] ), .B(\mem[41][5] ), .C(\mem[42][5] ), .D(
        \mem[43][5] ), .S0(n814), .S1(n838), .Y(n128) );
  MXI4X1 U823 ( .A(n80), .B(n78), .C(n79), .D(n77), .S0(n848), .S1(n844), .Y(
        n747) );
  MX4X1 U824 ( .A(\mem[108][6] ), .B(\mem[109][6] ), .C(\mem[110][6] ), .D(
        \mem[111][6] ), .S0(n811), .S1(n829), .Y(n77) );
  MX4X1 U825 ( .A(\mem[100][6] ), .B(\mem[101][6] ), .C(\mem[102][6] ), .D(
        \mem[103][6] ), .S0(n811), .S1(n838), .Y(n79) );
  MX4X1 U826 ( .A(\mem[104][6] ), .B(\mem[105][6] ), .C(\mem[106][6] ), .D(
        \mem[107][6] ), .S0(n811), .S1(n828), .Y(n78) );
  MXI4X1 U827 ( .A(n96), .B(n94), .C(n95), .D(n93), .S0(N29), .S1(n844), .Y(
        n751) );
  MX4X1 U828 ( .A(\mem[44][6] ), .B(\mem[45][6] ), .C(\mem[46][6] ), .D(
        \mem[47][6] ), .S0(n812), .S1(n835), .Y(n93) );
  MX4X1 U829 ( .A(\mem[36][6] ), .B(\mem[37][6] ), .C(\mem[38][6] ), .D(
        \mem[39][6] ), .S0(n812), .S1(n835), .Y(n95) );
  MX4X1 U830 ( .A(\mem[40][6] ), .B(\mem[41][6] ), .C(\mem[42][6] ), .D(
        \mem[43][6] ), .S0(n812), .S1(n835), .Y(n94) );
  MXI4X1 U831 ( .A(n46), .B(n44), .C(n45), .D(n43), .S0(n849), .S1(n844), .Y(
        n739) );
  MX4X1 U832 ( .A(\mem[108][7] ), .B(\mem[109][7] ), .C(\mem[110][7] ), .D(
        \mem[111][7] ), .S0(n808), .S1(n832), .Y(n43) );
  MX4X1 U833 ( .A(\mem[100][7] ), .B(\mem[101][7] ), .C(\mem[102][7] ), .D(
        \mem[103][7] ), .S0(n808), .S1(n832), .Y(n45) );
  MX4X1 U834 ( .A(\mem[104][7] ), .B(\mem[105][7] ), .C(\mem[106][7] ), .D(
        \mem[107][7] ), .S0(n808), .S1(n832), .Y(n44) );
  MXI4X1 U835 ( .A(n62), .B(n60), .C(n61), .D(n59), .S0(n848), .S1(n846), .Y(
        n743) );
  MX4X1 U836 ( .A(\mem[44][7] ), .B(\mem[45][7] ), .C(\mem[46][7] ), .D(
        \mem[47][7] ), .S0(n809), .S1(n833), .Y(n59) );
  MX4X1 U837 ( .A(\mem[36][7] ), .B(\mem[37][7] ), .C(\mem[38][7] ), .D(
        \mem[39][7] ), .S0(n810), .S1(n834), .Y(n61) );
  MX4X1 U838 ( .A(\mem[40][7] ), .B(\mem[41][7] ), .C(\mem[42][7] ), .D(
        \mem[43][7] ), .S0(n809), .S1(n833), .Y(n60) );
  MXI4X1 U839 ( .A(n12), .B(n10), .C(n11), .D(n9), .S0(n849), .S1(n844), .Y(
        n731) );
  MX4X1 U840 ( .A(valid_mem[108]), .B(valid_mem[109]), .C(valid_mem[110]), .D(
        valid_mem[111]), .S0(n806), .S1(n829), .Y(n9) );
  MX4X1 U841 ( .A(valid_mem[100]), .B(valid_mem[101]), .C(valid_mem[102]), .D(
        valid_mem[103]), .S0(n806), .S1(n835), .Y(n11) );
  MX4X1 U842 ( .A(valid_mem[104]), .B(valid_mem[105]), .C(valid_mem[106]), .D(
        valid_mem[107]), .S0(n806), .S1(n829), .Y(n10) );
  MXI4X1 U843 ( .A(n28), .B(n26), .C(n27), .D(n25), .S0(n849), .S1(n844), .Y(
        n735) );
  MX4X1 U844 ( .A(valid_mem[44]), .B(valid_mem[45]), .C(valid_mem[46]), .D(
        valid_mem[47]), .S0(n807), .S1(n831), .Y(n25) );
  MX4X1 U845 ( .A(valid_mem[36]), .B(valid_mem[37]), .C(valid_mem[38]), .D(
        valid_mem[39]), .S0(n807), .S1(n831), .Y(n27) );
  MX4X1 U846 ( .A(valid_mem[40]), .B(valid_mem[41]), .C(valid_mem[42]), .D(
        valid_mem[43]), .S0(n807), .S1(n831), .Y(n26) );
  NAND2X1 U847 ( .A(n152), .B(n153), .Y(n448) );
  OAI21XL U848 ( .A0(n870), .A1(n155), .B0(valid_mem[127]), .Y(n153) );
  NAND2X1 U849 ( .A(n212), .B(n213), .Y(n469) );
  OAI21XL U850 ( .A0(n170), .A1(n868), .B0(valid_mem[106]), .Y(n213) );
  NAND2X1 U851 ( .A(n344), .B(n345), .Y(n533) );
  OAI21XL U852 ( .A0(n170), .A1(n860), .B0(valid_mem[42]), .Y(n345) );
  NAND2X1 U853 ( .A(n352), .B(n353), .Y(n537) );
  OAI21XL U854 ( .A0(n182), .A1(n860), .B0(valid_mem[38]), .Y(n353) );
  NAND2X1 U855 ( .A(n377), .B(n378), .Y(n549) );
  OAI21XL U856 ( .A0(n170), .A1(n858), .B0(valid_mem[26]), .Y(n378) );
  NAND2X1 U857 ( .A(n385), .B(n386), .Y(n553) );
  OAI21XL U858 ( .A0(n182), .A1(n858), .B0(valid_mem[22]), .Y(n386) );
  NAND2X1 U859 ( .A(n201), .B(n202), .Y(n464) );
  OAI21XL U860 ( .A0(n155), .A1(n868), .B0(valid_mem[111]), .Y(n202) );
  NAND2X1 U861 ( .A(n204), .B(n205), .Y(n465) );
  OAI21XL U862 ( .A0(n158), .A1(n868), .B0(valid_mem[110]), .Y(n205) );
  NAND2X1 U863 ( .A(n206), .B(n207), .Y(n466) );
  OAI21XL U864 ( .A0(n161), .A1(n868), .B0(valid_mem[109]), .Y(n207) );
  NAND2X1 U865 ( .A(n208), .B(n209), .Y(n467) );
  OAI21XL U866 ( .A0(n164), .A1(n868), .B0(valid_mem[108]), .Y(n209) );
  NAND2X1 U867 ( .A(n210), .B(n211), .Y(n468) );
  OAI21XL U868 ( .A0(n167), .A1(n868), .B0(valid_mem[107]), .Y(n211) );
  NAND2X1 U869 ( .A(n214), .B(n215), .Y(n470) );
  OAI21XL U870 ( .A0(n173), .A1(n868), .B0(valid_mem[105]), .Y(n215) );
  NAND2X1 U871 ( .A(n216), .B(n217), .Y(n471) );
  OAI21XL U872 ( .A0(n176), .A1(n868), .B0(valid_mem[104]), .Y(n217) );
  NAND2X1 U873 ( .A(n220), .B(n221), .Y(n473) );
  OAI21XL U874 ( .A0(n182), .A1(n868), .B0(valid_mem[102]), .Y(n221) );
  NAND2X1 U875 ( .A(n245), .B(n246), .Y(n485) );
  OAI21XL U876 ( .A0(n170), .A1(n866), .B0(valid_mem[90]), .Y(n246) );
  NAND2X1 U877 ( .A(n253), .B(n254), .Y(n489) );
  OAI21XL U878 ( .A0(n182), .A1(n866), .B0(valid_mem[86]), .Y(n254) );
  NAND2X1 U879 ( .A(n261), .B(n262), .Y(n493) );
  OAI21XL U880 ( .A0(n194), .A1(n866), .B0(valid_mem[82]), .Y(n262) );
  NAND2X1 U881 ( .A(n278), .B(n279), .Y(n501) );
  OAI21XL U882 ( .A0(n170), .A1(n864), .B0(valid_mem[74]), .Y(n279) );
  NAND2X1 U883 ( .A(n286), .B(n287), .Y(n505) );
  OAI21XL U884 ( .A0(n182), .A1(n864), .B0(valid_mem[70]), .Y(n287) );
  NAND2X1 U885 ( .A(n294), .B(n295), .Y(n509) );
  OAI21XL U886 ( .A0(n194), .A1(n864), .B0(valid_mem[66]), .Y(n295) );
  NAND2X1 U887 ( .A(n311), .B(n312), .Y(n517) );
  OAI21XL U888 ( .A0(n170), .A1(n862), .B0(valid_mem[58]), .Y(n312) );
  NAND2X1 U889 ( .A(n218), .B(n219), .Y(n472) );
  OAI21XL U890 ( .A0(n179), .A1(n868), .B0(valid_mem[103]), .Y(n219) );
  NAND2X1 U891 ( .A(n222), .B(n223), .Y(n474) );
  OAI21XL U892 ( .A0(n185), .A1(n868), .B0(valid_mem[101]), .Y(n223) );
  NAND2X1 U893 ( .A(n224), .B(n225), .Y(n475) );
  OAI21XL U894 ( .A0(n188), .A1(n868), .B0(valid_mem[100]), .Y(n225) );
  NAND2X1 U895 ( .A(n228), .B(n229), .Y(n477) );
  OAI21XL U896 ( .A0(n194), .A1(n868), .B0(valid_mem[98]), .Y(n229) );
  NAND2X1 U897 ( .A(n226), .B(n227), .Y(n476) );
  OAI21XL U898 ( .A0(n191), .A1(n868), .B0(valid_mem[99]), .Y(n227) );
  NAND2X1 U899 ( .A(n230), .B(n231), .Y(n478) );
  OAI21XL U900 ( .A0(n197), .A1(n868), .B0(valid_mem[97]), .Y(n231) );
  NAND2X1 U901 ( .A(n232), .B(n233), .Y(n479) );
  OAI21XL U902 ( .A0(n200), .A1(n868), .B0(valid_mem[96]), .Y(n233) );
  NAND2X1 U903 ( .A(n234), .B(n235), .Y(n480) );
  OAI21XL U904 ( .A0(n155), .A1(n866), .B0(valid_mem[95]), .Y(n235) );
  NAND2X1 U905 ( .A(n237), .B(n238), .Y(n481) );
  OAI21XL U906 ( .A0(n158), .A1(n866), .B0(valid_mem[94]), .Y(n238) );
  NAND2X1 U907 ( .A(n239), .B(n240), .Y(n482) );
  OAI21XL U908 ( .A0(n161), .A1(n866), .B0(valid_mem[93]), .Y(n240) );
  NAND2X1 U909 ( .A(n241), .B(n242), .Y(n483) );
  OAI21XL U910 ( .A0(n164), .A1(n866), .B0(valid_mem[92]), .Y(n242) );
  NAND2X1 U911 ( .A(n243), .B(n244), .Y(n484) );
  OAI21XL U912 ( .A0(n167), .A1(n866), .B0(valid_mem[91]), .Y(n244) );
  NAND2X1 U913 ( .A(n247), .B(n248), .Y(n486) );
  OAI21XL U914 ( .A0(n173), .A1(n866), .B0(valid_mem[89]), .Y(n248) );
  NAND2X1 U915 ( .A(n249), .B(n250), .Y(n487) );
  OAI21XL U916 ( .A0(n176), .A1(n866), .B0(valid_mem[88]), .Y(n250) );
  NAND2X1 U917 ( .A(n251), .B(n252), .Y(n488) );
  OAI21XL U918 ( .A0(n179), .A1(n866), .B0(valid_mem[87]), .Y(n252) );
  NAND2X1 U919 ( .A(n255), .B(n256), .Y(n490) );
  OAI21XL U920 ( .A0(n185), .A1(n866), .B0(valid_mem[85]), .Y(n256) );
  NAND2X1 U921 ( .A(n257), .B(n258), .Y(n491) );
  OAI21XL U922 ( .A0(n188), .A1(n866), .B0(valid_mem[84]), .Y(n258) );
  NAND2X1 U923 ( .A(n259), .B(n260), .Y(n492) );
  OAI21XL U924 ( .A0(n191), .A1(n866), .B0(valid_mem[83]), .Y(n260) );
  NAND2X1 U925 ( .A(n263), .B(n264), .Y(n494) );
  OAI21XL U926 ( .A0(n197), .A1(n866), .B0(valid_mem[81]), .Y(n264) );
  NAND2X1 U927 ( .A(n265), .B(n266), .Y(n495) );
  OAI21XL U928 ( .A0(n200), .A1(n866), .B0(valid_mem[80]), .Y(n266) );
  NAND2X1 U929 ( .A(n267), .B(n268), .Y(n496) );
  OAI21XL U930 ( .A0(n155), .A1(n864), .B0(valid_mem[79]), .Y(n268) );
  NAND2X1 U931 ( .A(n270), .B(n271), .Y(n497) );
  OAI21XL U932 ( .A0(n158), .A1(n864), .B0(valid_mem[78]), .Y(n271) );
  NAND2X1 U933 ( .A(n272), .B(n273), .Y(n498) );
  OAI21XL U934 ( .A0(n161), .A1(n864), .B0(valid_mem[77]), .Y(n273) );
  NAND2X1 U935 ( .A(n274), .B(n275), .Y(n499) );
  OAI21XL U936 ( .A0(n164), .A1(n864), .B0(valid_mem[76]), .Y(n275) );
  NAND2X1 U937 ( .A(n276), .B(n277), .Y(n500) );
  OAI21XL U938 ( .A0(n167), .A1(n864), .B0(valid_mem[75]), .Y(n277) );
  NAND2X1 U939 ( .A(n280), .B(n281), .Y(n502) );
  OAI21XL U940 ( .A0(n173), .A1(n864), .B0(valid_mem[73]), .Y(n281) );
  NAND2X1 U941 ( .A(n282), .B(n283), .Y(n503) );
  OAI21XL U942 ( .A0(n176), .A1(n864), .B0(valid_mem[72]), .Y(n283) );
  NAND2X1 U943 ( .A(n284), .B(n285), .Y(n504) );
  OAI21XL U944 ( .A0(n179), .A1(n864), .B0(valid_mem[71]), .Y(n285) );
  NAND2X1 U945 ( .A(n288), .B(n289), .Y(n506) );
  OAI21XL U946 ( .A0(n185), .A1(n864), .B0(valid_mem[69]), .Y(n289) );
  NAND2X1 U947 ( .A(n290), .B(n291), .Y(n507) );
  OAI21XL U948 ( .A0(n188), .A1(n864), .B0(valid_mem[68]), .Y(n291) );
  NAND2X1 U949 ( .A(n292), .B(n293), .Y(n508) );
  OAI21XL U950 ( .A0(n191), .A1(n864), .B0(valid_mem[67]), .Y(n293) );
  NAND2X1 U951 ( .A(n296), .B(n297), .Y(n510) );
  OAI21XL U952 ( .A0(n197), .A1(n864), .B0(valid_mem[65]), .Y(n297) );
  NAND2X1 U953 ( .A(n298), .B(n299), .Y(n511) );
  OAI21XL U954 ( .A0(n200), .A1(n864), .B0(valid_mem[64]), .Y(n299) );
  NAND2X1 U955 ( .A(n300), .B(n301), .Y(n512) );
  OAI21XL U956 ( .A0(n155), .A1(n862), .B0(valid_mem[63]), .Y(n301) );
  NAND2X1 U957 ( .A(n303), .B(n304), .Y(n513) );
  OAI21XL U958 ( .A0(n158), .A1(n862), .B0(valid_mem[62]), .Y(n304) );
  NAND2X1 U959 ( .A(n305), .B(n306), .Y(n514) );
  OAI21XL U960 ( .A0(n161), .A1(n862), .B0(valid_mem[61]), .Y(n306) );
  NAND2X1 U961 ( .A(n307), .B(n308), .Y(n515) );
  OAI21XL U962 ( .A0(n164), .A1(n862), .B0(valid_mem[60]), .Y(n308) );
  NAND2X1 U963 ( .A(n309), .B(n310), .Y(n516) );
  OAI21XL U964 ( .A0(n167), .A1(n862), .B0(valid_mem[59]), .Y(n310) );
  NAND2X1 U965 ( .A(n313), .B(n314), .Y(n518) );
  OAI21XL U966 ( .A0(n173), .A1(n862), .B0(valid_mem[57]), .Y(n314) );
  NAND2X1 U967 ( .A(n315), .B(n316), .Y(n519) );
  OAI21XL U968 ( .A0(n176), .A1(n862), .B0(valid_mem[56]), .Y(n316) );
  NAND2X1 U969 ( .A(n319), .B(n320), .Y(n521) );
  OAI21XL U970 ( .A0(n182), .A1(n862), .B0(valid_mem[54]), .Y(n320) );
  NAND2X1 U971 ( .A(n317), .B(n318), .Y(n520) );
  OAI21XL U972 ( .A0(n179), .A1(n862), .B0(valid_mem[55]), .Y(n318) );
  NAND2X1 U973 ( .A(n321), .B(n322), .Y(n522) );
  OAI21XL U974 ( .A0(n185), .A1(n862), .B0(valid_mem[53]), .Y(n322) );
  NAND2X1 U975 ( .A(n323), .B(n324), .Y(n523) );
  OAI21XL U976 ( .A0(n188), .A1(n862), .B0(valid_mem[52]), .Y(n324) );
  NAND2X1 U977 ( .A(n327), .B(n328), .Y(n525) );
  OAI21XL U978 ( .A0(n194), .A1(n862), .B0(valid_mem[50]), .Y(n328) );
  NAND2X1 U979 ( .A(n325), .B(n326), .Y(n524) );
  OAI21XL U980 ( .A0(n191), .A1(n862), .B0(valid_mem[51]), .Y(n326) );
  NAND2X1 U981 ( .A(n329), .B(n330), .Y(n526) );
  OAI21XL U982 ( .A0(n197), .A1(n862), .B0(valid_mem[49]), .Y(n330) );
  NAND2X1 U983 ( .A(n331), .B(n332), .Y(n527) );
  OAI21XL U984 ( .A0(n200), .A1(n862), .B0(valid_mem[48]), .Y(n332) );
  NAND2X1 U985 ( .A(n333), .B(n334), .Y(n528) );
  OAI21XL U986 ( .A0(n155), .A1(n860), .B0(valid_mem[47]), .Y(n334) );
  NAND2X1 U987 ( .A(n336), .B(n337), .Y(n529) );
  OAI21XL U988 ( .A0(n158), .A1(n860), .B0(valid_mem[46]), .Y(n337) );
  NAND2X1 U989 ( .A(n338), .B(n339), .Y(n530) );
  OAI21XL U990 ( .A0(n161), .A1(n860), .B0(valid_mem[45]), .Y(n339) );
  NAND2X1 U991 ( .A(n340), .B(n341), .Y(n531) );
  OAI21XL U992 ( .A0(n164), .A1(n860), .B0(valid_mem[44]), .Y(n341) );
  NAND2X1 U993 ( .A(n342), .B(n343), .Y(n532) );
  OAI21XL U994 ( .A0(n167), .A1(n860), .B0(valid_mem[43]), .Y(n343) );
  NAND2X1 U995 ( .A(n346), .B(n347), .Y(n534) );
  OAI21XL U996 ( .A0(n173), .A1(n860), .B0(valid_mem[41]), .Y(n347) );
  NAND2X1 U997 ( .A(n348), .B(n349), .Y(n535) );
  OAI21XL U998 ( .A0(n176), .A1(n860), .B0(valid_mem[40]), .Y(n349) );
  NAND2X1 U999 ( .A(n350), .B(n351), .Y(n536) );
  OAI21XL U1000 ( .A0(n179), .A1(n860), .B0(valid_mem[39]), .Y(n351) );
  NAND2X1 U1001 ( .A(n354), .B(n355), .Y(n538) );
  OAI21XL U1002 ( .A0(n185), .A1(n860), .B0(valid_mem[37]), .Y(n355) );
  NAND2X1 U1003 ( .A(n356), .B(n357), .Y(n539) );
  OAI21XL U1004 ( .A0(n188), .A1(n860), .B0(valid_mem[36]), .Y(n357) );
  NAND2X1 U1005 ( .A(n360), .B(n361), .Y(n541) );
  OAI21XL U1006 ( .A0(n194), .A1(n860), .B0(valid_mem[34]), .Y(n361) );
  NAND2X1 U1007 ( .A(n358), .B(n359), .Y(n540) );
  OAI21XL U1008 ( .A0(n191), .A1(n860), .B0(valid_mem[35]), .Y(n359) );
  NAND2X1 U1009 ( .A(n362), .B(n363), .Y(n542) );
  OAI21XL U1010 ( .A0(n197), .A1(n860), .B0(valid_mem[33]), .Y(n363) );
  NAND2X1 U1011 ( .A(n364), .B(n365), .Y(n543) );
  OAI21XL U1012 ( .A0(n200), .A1(n860), .B0(valid_mem[32]), .Y(n365) );
  NAND2X1 U1013 ( .A(n366), .B(n367), .Y(n544) );
  OAI21XL U1014 ( .A0(n155), .A1(n858), .B0(valid_mem[31]), .Y(n367) );
  NAND2X1 U1015 ( .A(n369), .B(n370), .Y(n545) );
  OAI21XL U1016 ( .A0(n158), .A1(n858), .B0(valid_mem[30]), .Y(n370) );
  NAND2X1 U1017 ( .A(n371), .B(n372), .Y(n546) );
  OAI21XL U1018 ( .A0(n161), .A1(n858), .B0(valid_mem[29]), .Y(n372) );
  NAND2X1 U1019 ( .A(n373), .B(n374), .Y(n547) );
  OAI21XL U1020 ( .A0(n164), .A1(n858), .B0(valid_mem[28]), .Y(n374) );
  NAND2X1 U1021 ( .A(n375), .B(n376), .Y(n548) );
  OAI21XL U1022 ( .A0(n167), .A1(n858), .B0(valid_mem[27]), .Y(n376) );
  NAND2X1 U1023 ( .A(n379), .B(n380), .Y(n550) );
  OAI21XL U1024 ( .A0(n173), .A1(n858), .B0(valid_mem[25]), .Y(n380) );
  NAND2X1 U1025 ( .A(n381), .B(n382), .Y(n551) );
  OAI21XL U1026 ( .A0(n176), .A1(n858), .B0(valid_mem[24]), .Y(n382) );
  NAND2X1 U1027 ( .A(n383), .B(n384), .Y(n552) );
  OAI21XL U1028 ( .A0(n179), .A1(n858), .B0(valid_mem[23]), .Y(n384) );
  NAND2X1 U1029 ( .A(n387), .B(n388), .Y(n554) );
  OAI21XL U1030 ( .A0(n185), .A1(n858), .B0(valid_mem[21]), .Y(n388) );
  NAND2X1 U1031 ( .A(n389), .B(n390), .Y(n555) );
  OAI21XL U1032 ( .A0(n188), .A1(n858), .B0(valid_mem[20]), .Y(n390) );
  NAND2X1 U1033 ( .A(n393), .B(n394), .Y(n557) );
  OAI21XL U1034 ( .A0(n194), .A1(n858), .B0(valid_mem[18]), .Y(n394) );
  NAND2X1 U1035 ( .A(n391), .B(n392), .Y(n556) );
  OAI21XL U1036 ( .A0(n191), .A1(n858), .B0(valid_mem[19]), .Y(n392) );
  NAND2X1 U1037 ( .A(n395), .B(n396), .Y(n558) );
  OAI21XL U1038 ( .A0(n197), .A1(n858), .B0(valid_mem[17]), .Y(n396) );
  NAND2X1 U1039 ( .A(n397), .B(n398), .Y(n559) );
  OAI21XL U1040 ( .A0(n200), .A1(n858), .B0(valid_mem[16]), .Y(n398) );
  NAND2X1 U1041 ( .A(n410), .B(n411), .Y(n565) );
  OAI21XL U1042 ( .A0(n170), .A1(n856), .B0(valid_mem[10]), .Y(n411) );
  NAND2X1 U1043 ( .A(n399), .B(n400), .Y(n560) );
  OAI21XL U1044 ( .A0(n155), .A1(n856), .B0(valid_mem[15]), .Y(n400) );
  NAND2X1 U1045 ( .A(n402), .B(n403), .Y(n561) );
  OAI21XL U1046 ( .A0(n158), .A1(n856), .B0(valid_mem[14]), .Y(n403) );
  NAND2X1 U1047 ( .A(n404), .B(n405), .Y(n562) );
  OAI21XL U1048 ( .A0(n161), .A1(n856), .B0(valid_mem[13]), .Y(n405) );
  NAND2X1 U1049 ( .A(n406), .B(n407), .Y(n563) );
  OAI21XL U1050 ( .A0(n164), .A1(n856), .B0(valid_mem[12]), .Y(n407) );
  NAND2X1 U1051 ( .A(n408), .B(n409), .Y(n564) );
  OAI21XL U1052 ( .A0(n167), .A1(n856), .B0(valid_mem[11]), .Y(n409) );
  NAND2X1 U1053 ( .A(n412), .B(n413), .Y(n566) );
  OAI21XL U1054 ( .A0(n173), .A1(n856), .B0(valid_mem[9]), .Y(n413) );
  NAND2X1 U1055 ( .A(n414), .B(n415), .Y(n567) );
  OAI21XL U1056 ( .A0(n176), .A1(n856), .B0(valid_mem[8]), .Y(n415) );
  NAND2X1 U1057 ( .A(n418), .B(n419), .Y(n569) );
  OAI21XL U1058 ( .A0(n182), .A1(n856), .B0(valid_mem[6]), .Y(n419) );
  NAND2X1 U1059 ( .A(n416), .B(n417), .Y(n568) );
  OAI21XL U1060 ( .A0(n179), .A1(n856), .B0(valid_mem[7]), .Y(n417) );
  NAND2X1 U1061 ( .A(n420), .B(n421), .Y(n570) );
  OAI21XL U1062 ( .A0(n185), .A1(n856), .B0(valid_mem[5]), .Y(n421) );
  NAND2X1 U1063 ( .A(n422), .B(n423), .Y(n571) );
  OAI21XL U1064 ( .A0(n188), .A1(n856), .B0(valid_mem[4]), .Y(n423) );
  NAND2X1 U1065 ( .A(n426), .B(n427), .Y(n573) );
  OAI21XL U1066 ( .A0(n194), .A1(n856), .B0(valid_mem[2]), .Y(n427) );
  NAND2X1 U1067 ( .A(n424), .B(n425), .Y(n572) );
  OAI21XL U1068 ( .A0(n191), .A1(n856), .B0(valid_mem[3]), .Y(n425) );
  NAND2X1 U1069 ( .A(n428), .B(n429), .Y(n574) );
  OAI21XL U1070 ( .A0(n197), .A1(n856), .B0(valid_mem[1]), .Y(n429) );
  NAND2X1 U1071 ( .A(n430), .B(n431), .Y(n575) );
  OAI21XL U1072 ( .A0(n200), .A1(n856), .B0(valid_mem[0]), .Y(n431) );
endmodule


module up_counter_WIDTH7_0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module up_counter_WIDTH7_0 ( clk, rst, en, clr, count );
  output [6:0] count;
  input clk, rst, en, clr;
  wire   n18, N4, N5, N6, N7, N8, N9, N10, n1, n2, n4, n11, n12, n13, n14, n15,
         n16, n17;

  up_counter_WIDTH7_0_DW01_inc_0 add_18 ( .A({count[6], n18, count[4:0]}), 
        .SUM({N10, N9, N8, N7, N6, N5, N4}) );
  DFFRX1 \count_reg[5]  ( .D(n16), .CK(clk), .RN(n11), .Q(n18), .QN(n2) );
  DFFRX1 \count_reg[3]  ( .D(n14), .CK(clk), .RN(n11), .Q(count[3]) );
  DFFRX1 \count_reg[2]  ( .D(n13), .CK(clk), .RN(n11), .Q(count[2]) );
  DFFRX1 \count_reg[1]  ( .D(n12), .CK(clk), .RN(n11), .Q(count[1]) );
  DFFRX2 \count_reg[6]  ( .D(n17), .CK(clk), .RN(n11), .Q(count[6]) );
  DFFRX2 \count_reg[0]  ( .D(n1), .CK(clk), .RN(n11), .Q(count[0]) );
  DFFRX2 \count_reg[4]  ( .D(n15), .CK(clk), .RN(n11), .Q(count[4]) );
  AO22X1 U3 ( .A0(N4), .A1(en), .B0(count[0]), .B1(n4), .Y(n1) );
  CLKINVX1 U4 ( .A(n2), .Y(count[5]) );
  CLKINVX1 U5 ( .A(en), .Y(n4) );
  INVX3 U6 ( .A(rst), .Y(n11) );
  AO22X1 U7 ( .A0(count[6]), .A1(n4), .B0(N10), .B1(en), .Y(n17) );
  AO22XL U8 ( .A0(count[4]), .A1(n4), .B0(N8), .B1(en), .Y(n15) );
  AO22XL U9 ( .A0(n18), .A1(n4), .B0(N9), .B1(en), .Y(n16) );
  AO22X1 U10 ( .A0(count[3]), .A1(n4), .B0(N7), .B1(en), .Y(n14) );
  AO22X1 U11 ( .A0(count[1]), .A1(n4), .B0(N5), .B1(en), .Y(n12) );
  AO22X1 U12 ( .A0(count[2]), .A1(n4), .B0(N6), .B1(en), .Y(n13) );
endmodule


module line_buffer_0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module line_buffer_0 ( clk, rst, en, data_in, data_out, valid );
  input [7:0] data_in;
  output [7:0] data_out;
  input clk, rst, en;
  output valid;
  wire   N26, N27, N28, N29, N30, N31, N32, \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] ,
         \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] ,
         \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] ,
         \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] ,
         \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] ,
         \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[15][7] , \mem[15][6] ,
         \mem[15][5] , \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] ,
         \mem[15][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] , \mem[16][4] ,
         \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] ,
         \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] ,
         \mem[19][7] , \mem[19][6] , \mem[19][5] , \mem[19][4] , \mem[19][3] ,
         \mem[19][2] , \mem[19][1] , \mem[19][0] , \mem[20][7] , \mem[20][6] ,
         \mem[20][5] , \mem[20][4] , \mem[20][3] , \mem[20][2] , \mem[20][1] ,
         \mem[20][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] , \mem[21][4] ,
         \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] ,
         \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] ,
         \mem[24][7] , \mem[24][6] , \mem[24][5] , \mem[24][4] , \mem[24][3] ,
         \mem[24][2] , \mem[24][1] , \mem[24][0] , \mem[25][7] , \mem[25][6] ,
         \mem[25][5] , \mem[25][4] , \mem[25][3] , \mem[25][2] , \mem[25][1] ,
         \mem[25][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] , \mem[26][4] ,
         \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] ,
         \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] ,
         \mem[29][7] , \mem[29][6] , \mem[29][5] , \mem[29][4] , \mem[29][3] ,
         \mem[29][2] , \mem[29][1] , \mem[29][0] , \mem[30][7] , \mem[30][6] ,
         \mem[30][5] , \mem[30][4] , \mem[30][3] , \mem[30][2] , \mem[30][1] ,
         \mem[30][0] , \mem[31][7] , \mem[31][6] , \mem[31][5] , \mem[31][4] ,
         \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] , \mem[32][7] ,
         \mem[32][6] , \mem[32][5] , \mem[32][4] , \mem[32][3] , \mem[32][2] ,
         \mem[32][1] , \mem[32][0] , \mem[33][7] , \mem[33][6] , \mem[33][5] ,
         \mem[33][4] , \mem[33][3] , \mem[33][2] , \mem[33][1] , \mem[33][0] ,
         \mem[34][7] , \mem[34][6] , \mem[34][5] , \mem[34][4] , \mem[34][3] ,
         \mem[34][2] , \mem[34][1] , \mem[34][0] , \mem[35][7] , \mem[35][6] ,
         \mem[35][5] , \mem[35][4] , \mem[35][3] , \mem[35][2] , \mem[35][1] ,
         \mem[35][0] , \mem[36][7] , \mem[36][6] , \mem[36][5] , \mem[36][4] ,
         \mem[36][3] , \mem[36][2] , \mem[36][1] , \mem[36][0] , \mem[37][7] ,
         \mem[37][6] , \mem[37][5] , \mem[37][4] , \mem[37][3] , \mem[37][2] ,
         \mem[37][1] , \mem[37][0] , \mem[38][7] , \mem[38][6] , \mem[38][5] ,
         \mem[38][4] , \mem[38][3] , \mem[38][2] , \mem[38][1] , \mem[38][0] ,
         \mem[39][7] , \mem[39][6] , \mem[39][5] , \mem[39][4] , \mem[39][3] ,
         \mem[39][2] , \mem[39][1] , \mem[39][0] , \mem[40][7] , \mem[40][6] ,
         \mem[40][5] , \mem[40][4] , \mem[40][3] , \mem[40][2] , \mem[40][1] ,
         \mem[40][0] , \mem[41][7] , \mem[41][6] , \mem[41][5] , \mem[41][4] ,
         \mem[41][3] , \mem[41][2] , \mem[41][1] , \mem[41][0] , \mem[42][7] ,
         \mem[42][6] , \mem[42][5] , \mem[42][4] , \mem[42][3] , \mem[42][2] ,
         \mem[42][1] , \mem[42][0] , \mem[43][7] , \mem[43][6] , \mem[43][5] ,
         \mem[43][4] , \mem[43][3] , \mem[43][2] , \mem[43][1] , \mem[43][0] ,
         \mem[44][7] , \mem[44][6] , \mem[44][5] , \mem[44][4] , \mem[44][3] ,
         \mem[44][2] , \mem[44][1] , \mem[44][0] , \mem[45][7] , \mem[45][6] ,
         \mem[45][5] , \mem[45][4] , \mem[45][3] , \mem[45][2] , \mem[45][1] ,
         \mem[45][0] , \mem[46][7] , \mem[46][6] , \mem[46][5] , \mem[46][4] ,
         \mem[46][3] , \mem[46][2] , \mem[46][1] , \mem[46][0] , \mem[47][7] ,
         \mem[47][6] , \mem[47][5] , \mem[47][4] , \mem[47][3] , \mem[47][2] ,
         \mem[47][1] , \mem[47][0] , \mem[48][7] , \mem[48][6] , \mem[48][5] ,
         \mem[48][4] , \mem[48][3] , \mem[48][2] , \mem[48][1] , \mem[48][0] ,
         \mem[49][7] , \mem[49][6] , \mem[49][5] , \mem[49][4] , \mem[49][3] ,
         \mem[49][2] , \mem[49][1] , \mem[49][0] , \mem[50][7] , \mem[50][6] ,
         \mem[50][5] , \mem[50][4] , \mem[50][3] , \mem[50][2] , \mem[50][1] ,
         \mem[50][0] , \mem[51][7] , \mem[51][6] , \mem[51][5] , \mem[51][4] ,
         \mem[51][3] , \mem[51][2] , \mem[51][1] , \mem[51][0] , \mem[52][7] ,
         \mem[52][6] , \mem[52][5] , \mem[52][4] , \mem[52][3] , \mem[52][2] ,
         \mem[52][1] , \mem[52][0] , \mem[53][7] , \mem[53][6] , \mem[53][5] ,
         \mem[53][4] , \mem[53][3] , \mem[53][2] , \mem[53][1] , \mem[53][0] ,
         \mem[54][7] , \mem[54][6] , \mem[54][5] , \mem[54][4] , \mem[54][3] ,
         \mem[54][2] , \mem[54][1] , \mem[54][0] , \mem[55][7] , \mem[55][6] ,
         \mem[55][5] , \mem[55][4] , \mem[55][3] , \mem[55][2] , \mem[55][1] ,
         \mem[55][0] , \mem[56][7] , \mem[56][6] , \mem[56][5] , \mem[56][4] ,
         \mem[56][3] , \mem[56][2] , \mem[56][1] , \mem[56][0] , \mem[57][7] ,
         \mem[57][6] , \mem[57][5] , \mem[57][4] , \mem[57][3] , \mem[57][2] ,
         \mem[57][1] , \mem[57][0] , \mem[58][7] , \mem[58][6] , \mem[58][5] ,
         \mem[58][4] , \mem[58][3] , \mem[58][2] , \mem[58][1] , \mem[58][0] ,
         \mem[59][7] , \mem[59][6] , \mem[59][5] , \mem[59][4] , \mem[59][3] ,
         \mem[59][2] , \mem[59][1] , \mem[59][0] , \mem[60][7] , \mem[60][6] ,
         \mem[60][5] , \mem[60][4] , \mem[60][3] , \mem[60][2] , \mem[60][1] ,
         \mem[60][0] , \mem[61][7] , \mem[61][6] , \mem[61][5] , \mem[61][4] ,
         \mem[61][3] , \mem[61][2] , \mem[61][1] , \mem[61][0] , \mem[62][7] ,
         \mem[62][6] , \mem[62][5] , \mem[62][4] , \mem[62][3] , \mem[62][2] ,
         \mem[62][1] , \mem[62][0] , \mem[63][7] , \mem[63][6] , \mem[63][5] ,
         \mem[63][4] , \mem[63][3] , \mem[63][2] , \mem[63][1] , \mem[63][0] ,
         \mem[64][7] , \mem[64][6] , \mem[64][5] , \mem[64][4] , \mem[64][3] ,
         \mem[64][2] , \mem[64][1] , \mem[64][0] , \mem[65][7] , \mem[65][6] ,
         \mem[65][5] , \mem[65][4] , \mem[65][3] , \mem[65][2] , \mem[65][1] ,
         \mem[65][0] , \mem[66][7] , \mem[66][6] , \mem[66][5] , \mem[66][4] ,
         \mem[66][3] , \mem[66][2] , \mem[66][1] , \mem[66][0] , \mem[67][7] ,
         \mem[67][6] , \mem[67][5] , \mem[67][4] , \mem[67][3] , \mem[67][2] ,
         \mem[67][1] , \mem[67][0] , \mem[68][7] , \mem[68][6] , \mem[68][5] ,
         \mem[68][4] , \mem[68][3] , \mem[68][2] , \mem[68][1] , \mem[68][0] ,
         \mem[69][7] , \mem[69][6] , \mem[69][5] , \mem[69][4] , \mem[69][3] ,
         \mem[69][2] , \mem[69][1] , \mem[69][0] , \mem[70][7] , \mem[70][6] ,
         \mem[70][5] , \mem[70][4] , \mem[70][3] , \mem[70][2] , \mem[70][1] ,
         \mem[70][0] , \mem[71][7] , \mem[71][6] , \mem[71][5] , \mem[71][4] ,
         \mem[71][3] , \mem[71][2] , \mem[71][1] , \mem[71][0] , \mem[72][7] ,
         \mem[72][6] , \mem[72][5] , \mem[72][4] , \mem[72][3] , \mem[72][2] ,
         \mem[72][1] , \mem[72][0] , \mem[73][7] , \mem[73][6] , \mem[73][5] ,
         \mem[73][4] , \mem[73][3] , \mem[73][2] , \mem[73][1] , \mem[73][0] ,
         \mem[74][7] , \mem[74][6] , \mem[74][5] , \mem[74][4] , \mem[74][3] ,
         \mem[74][2] , \mem[74][1] , \mem[74][0] , \mem[75][7] , \mem[75][6] ,
         \mem[75][5] , \mem[75][4] , \mem[75][3] , \mem[75][2] , \mem[75][1] ,
         \mem[75][0] , \mem[76][7] , \mem[76][6] , \mem[76][5] , \mem[76][4] ,
         \mem[76][3] , \mem[76][2] , \mem[76][1] , \mem[76][0] , \mem[77][7] ,
         \mem[77][6] , \mem[77][5] , \mem[77][4] , \mem[77][3] , \mem[77][2] ,
         \mem[77][1] , \mem[77][0] , \mem[78][7] , \mem[78][6] , \mem[78][5] ,
         \mem[78][4] , \mem[78][3] , \mem[78][2] , \mem[78][1] , \mem[78][0] ,
         \mem[79][7] , \mem[79][6] , \mem[79][5] , \mem[79][4] , \mem[79][3] ,
         \mem[79][2] , \mem[79][1] , \mem[79][0] , \mem[80][7] , \mem[80][6] ,
         \mem[80][5] , \mem[80][4] , \mem[80][3] , \mem[80][2] , \mem[80][1] ,
         \mem[80][0] , \mem[81][7] , \mem[81][6] , \mem[81][5] , \mem[81][4] ,
         \mem[81][3] , \mem[81][2] , \mem[81][1] , \mem[81][0] , \mem[82][7] ,
         \mem[82][6] , \mem[82][5] , \mem[82][4] , \mem[82][3] , \mem[82][2] ,
         \mem[82][1] , \mem[82][0] , \mem[83][7] , \mem[83][6] , \mem[83][5] ,
         \mem[83][4] , \mem[83][3] , \mem[83][2] , \mem[83][1] , \mem[83][0] ,
         \mem[84][7] , \mem[84][6] , \mem[84][5] , \mem[84][4] , \mem[84][3] ,
         \mem[84][2] , \mem[84][1] , \mem[84][0] , \mem[85][7] , \mem[85][6] ,
         \mem[85][5] , \mem[85][4] , \mem[85][3] , \mem[85][2] , \mem[85][1] ,
         \mem[85][0] , \mem[86][7] , \mem[86][6] , \mem[86][5] , \mem[86][4] ,
         \mem[86][3] , \mem[86][2] , \mem[86][1] , \mem[86][0] , \mem[87][7] ,
         \mem[87][6] , \mem[87][5] , \mem[87][4] , \mem[87][3] , \mem[87][2] ,
         \mem[87][1] , \mem[87][0] , \mem[88][7] , \mem[88][6] , \mem[88][5] ,
         \mem[88][4] , \mem[88][3] , \mem[88][2] , \mem[88][1] , \mem[88][0] ,
         \mem[89][7] , \mem[89][6] , \mem[89][5] , \mem[89][4] , \mem[89][3] ,
         \mem[89][2] , \mem[89][1] , \mem[89][0] , \mem[90][7] , \mem[90][6] ,
         \mem[90][5] , \mem[90][4] , \mem[90][3] , \mem[90][2] , \mem[90][1] ,
         \mem[90][0] , \mem[91][7] , \mem[91][6] , \mem[91][5] , \mem[91][4] ,
         \mem[91][3] , \mem[91][2] , \mem[91][1] , \mem[91][0] , \mem[92][7] ,
         \mem[92][6] , \mem[92][5] , \mem[92][4] , \mem[92][3] , \mem[92][2] ,
         \mem[92][1] , \mem[92][0] , \mem[93][7] , \mem[93][6] , \mem[93][5] ,
         \mem[93][4] , \mem[93][3] , \mem[93][2] , \mem[93][1] , \mem[93][0] ,
         \mem[94][7] , \mem[94][6] , \mem[94][5] , \mem[94][4] , \mem[94][3] ,
         \mem[94][2] , \mem[94][1] , \mem[94][0] , \mem[95][7] , \mem[95][6] ,
         \mem[95][5] , \mem[95][4] , \mem[95][3] , \mem[95][2] , \mem[95][1] ,
         \mem[95][0] , \mem[96][7] , \mem[96][6] , \mem[96][5] , \mem[96][4] ,
         \mem[96][3] , \mem[96][2] , \mem[96][1] , \mem[96][0] , \mem[97][7] ,
         \mem[97][6] , \mem[97][5] , \mem[97][4] , \mem[97][3] , \mem[97][2] ,
         \mem[97][1] , \mem[97][0] , \mem[98][7] , \mem[98][6] , \mem[98][5] ,
         \mem[98][4] , \mem[98][3] , \mem[98][2] , \mem[98][1] , \mem[98][0] ,
         \mem[99][7] , \mem[99][6] , \mem[99][5] , \mem[99][4] , \mem[99][3] ,
         \mem[99][2] , \mem[99][1] , \mem[99][0] , \mem[100][7] ,
         \mem[100][6] , \mem[100][5] , \mem[100][4] , \mem[100][3] ,
         \mem[100][2] , \mem[100][1] , \mem[100][0] , \mem[101][7] ,
         \mem[101][6] , \mem[101][5] , \mem[101][4] , \mem[101][3] ,
         \mem[101][2] , \mem[101][1] , \mem[101][0] , \mem[102][7] ,
         \mem[102][6] , \mem[102][5] , \mem[102][4] , \mem[102][3] ,
         \mem[102][2] , \mem[102][1] , \mem[102][0] , \mem[103][7] ,
         \mem[103][6] , \mem[103][5] , \mem[103][4] , \mem[103][3] ,
         \mem[103][2] , \mem[103][1] , \mem[103][0] , \mem[104][7] ,
         \mem[104][6] , \mem[104][5] , \mem[104][4] , \mem[104][3] ,
         \mem[104][2] , \mem[104][1] , \mem[104][0] , \mem[105][7] ,
         \mem[105][6] , \mem[105][5] , \mem[105][4] , \mem[105][3] ,
         \mem[105][2] , \mem[105][1] , \mem[105][0] , \mem[106][7] ,
         \mem[106][6] , \mem[106][5] , \mem[106][4] , \mem[106][3] ,
         \mem[106][2] , \mem[106][1] , \mem[106][0] , \mem[107][7] ,
         \mem[107][6] , \mem[107][5] , \mem[107][4] , \mem[107][3] ,
         \mem[107][2] , \mem[107][1] , \mem[107][0] , \mem[108][7] ,
         \mem[108][6] , \mem[108][5] , \mem[108][4] , \mem[108][3] ,
         \mem[108][2] , \mem[108][1] , \mem[108][0] , \mem[109][7] ,
         \mem[109][6] , \mem[109][5] , \mem[109][4] , \mem[109][3] ,
         \mem[109][2] , \mem[109][1] , \mem[109][0] , \mem[110][7] ,
         \mem[110][6] , \mem[110][5] , \mem[110][4] , \mem[110][3] ,
         \mem[110][2] , \mem[110][1] , \mem[110][0] , \mem[111][7] ,
         \mem[111][6] , \mem[111][5] , \mem[111][4] , \mem[111][3] ,
         \mem[111][2] , \mem[111][1] , \mem[111][0] , \mem[112][7] ,
         \mem[112][6] , \mem[112][5] , \mem[112][4] , \mem[112][3] ,
         \mem[112][2] , \mem[112][1] , \mem[112][0] , \mem[113][7] ,
         \mem[113][6] , \mem[113][5] , \mem[113][4] , \mem[113][3] ,
         \mem[113][2] , \mem[113][1] , \mem[113][0] , \mem[114][7] ,
         \mem[114][6] , \mem[114][5] , \mem[114][4] , \mem[114][3] ,
         \mem[114][2] , \mem[114][1] , \mem[114][0] , \mem[115][7] ,
         \mem[115][6] , \mem[115][5] , \mem[115][4] , \mem[115][3] ,
         \mem[115][2] , \mem[115][1] , \mem[115][0] , \mem[116][7] ,
         \mem[116][6] , \mem[116][5] , \mem[116][4] , \mem[116][3] ,
         \mem[116][2] , \mem[116][1] , \mem[116][0] , \mem[117][7] ,
         \mem[117][6] , \mem[117][5] , \mem[117][4] , \mem[117][3] ,
         \mem[117][2] , \mem[117][1] , \mem[117][0] , \mem[118][7] ,
         \mem[118][6] , \mem[118][5] , \mem[118][4] , \mem[118][3] ,
         \mem[118][2] , \mem[118][1] , \mem[118][0] , \mem[119][7] ,
         \mem[119][6] , \mem[119][5] , \mem[119][4] , \mem[119][3] ,
         \mem[119][2] , \mem[119][1] , \mem[119][0] , \mem[120][7] ,
         \mem[120][6] , \mem[120][5] , \mem[120][4] , \mem[120][3] ,
         \mem[120][2] , \mem[120][1] , \mem[120][0] , \mem[121][7] ,
         \mem[121][6] , \mem[121][5] , \mem[121][4] , \mem[121][3] ,
         \mem[121][2] , \mem[121][1] , \mem[121][0] , \mem[122][7] ,
         \mem[122][6] , \mem[122][5] , \mem[122][4] , \mem[122][3] ,
         \mem[122][2] , \mem[122][1] , \mem[122][0] , \mem[123][7] ,
         \mem[123][6] , \mem[123][5] , \mem[123][4] , \mem[123][3] ,
         \mem[123][2] , \mem[123][1] , \mem[123][0] , \mem[124][7] ,
         \mem[124][6] , \mem[124][5] , \mem[124][4] , \mem[124][3] ,
         \mem[124][2] , \mem[124][1] , \mem[124][0] , \mem[125][7] ,
         \mem[125][6] , \mem[125][5] , \mem[125][4] , \mem[125][3] ,
         \mem[125][2] , \mem[125][1] , \mem[125][0] , \mem[126][7] ,
         \mem[126][6] , \mem[126][5] , \mem[126][4] , \mem[126][3] ,
         \mem[126][2] , \mem[126][1] , \mem[126][0] , \mem[127][7] ,
         \mem[127][6] , \mem[127][5] , \mem[127][4] , \mem[127][3] ,
         \mem[127][2] , \mem[127][1] , \mem[127][0] , N33, N34, N35, N36, N37,
         N38, N39, N40, N41, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n435,
         n436, n437, n438, n439, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488;
  wire   [6:0] write_counter_count;
  wire   [0:127] valid_mem;

  up_counter_WIDTH7_0 write_counter ( .clk(clk), .rst(rst), .en(n871), .clr(
        1'b0), .count(write_counter_count) );
  line_buffer_0_DW01_inc_0 add_15 ( .A(write_counter_count), .SUM({N32, N31, 
        N30, N29, N28, N27, N26}) );
  EDFFX1 \mem_reg[1][7]  ( .D(n915), .E(n963), .CK(clk), .Q(\mem[1][7] ) );
  EDFFX1 \mem_reg[1][6]  ( .D(n909), .E(n963), .CK(clk), .Q(\mem[1][6] ) );
  EDFFX1 \mem_reg[1][5]  ( .D(n903), .E(n963), .CK(clk), .Q(\mem[1][5] ) );
  EDFFX1 \mem_reg[1][4]  ( .D(n897), .E(n963), .CK(clk), .Q(\mem[1][4] ) );
  EDFFX1 \mem_reg[1][3]  ( .D(n891), .E(n963), .CK(clk), .Q(\mem[1][3] ) );
  EDFFX1 \mem_reg[1][2]  ( .D(n885), .E(n963), .CK(clk), .Q(\mem[1][2] ) );
  EDFFX1 \mem_reg[1][1]  ( .D(n879), .E(n963), .CK(clk), .Q(\mem[1][1] ) );
  EDFFX1 \mem_reg[1][0]  ( .D(n873), .E(n963), .CK(clk), .Q(\mem[1][0] ) );
  EDFFX1 \mem_reg[5][7]  ( .D(n914), .E(n972), .CK(clk), .Q(\mem[5][7] ) );
  EDFFX1 \mem_reg[5][6]  ( .D(n908), .E(n972), .CK(clk), .Q(\mem[5][6] ) );
  EDFFX1 \mem_reg[5][5]  ( .D(n902), .E(n972), .CK(clk), .Q(\mem[5][5] ) );
  EDFFX1 \mem_reg[5][4]  ( .D(n896), .E(n972), .CK(clk), .Q(\mem[5][4] ) );
  EDFFX1 \mem_reg[5][3]  ( .D(n890), .E(n972), .CK(clk), .Q(\mem[5][3] ) );
  EDFFX1 \mem_reg[5][2]  ( .D(n884), .E(n972), .CK(clk), .Q(\mem[5][2] ) );
  EDFFX1 \mem_reg[5][1]  ( .D(n878), .E(n972), .CK(clk), .Q(\mem[5][1] ) );
  EDFFX1 \mem_reg[5][0]  ( .D(n872), .E(n972), .CK(clk), .Q(\mem[5][0] ) );
  EDFFX1 \mem_reg[9][7]  ( .D(n919), .E(n981), .CK(clk), .Q(\mem[9][7] ) );
  EDFFX1 \mem_reg[9][6]  ( .D(n913), .E(n981), .CK(clk), .Q(\mem[9][6] ) );
  EDFFX1 \mem_reg[9][5]  ( .D(n907), .E(n981), .CK(clk), .Q(\mem[9][5] ) );
  EDFFX1 \mem_reg[9][4]  ( .D(n901), .E(n981), .CK(clk), .Q(\mem[9][4] ) );
  EDFFX1 \mem_reg[9][3]  ( .D(n895), .E(n981), .CK(clk), .Q(\mem[9][3] ) );
  EDFFX1 \mem_reg[9][2]  ( .D(n889), .E(n981), .CK(clk), .Q(\mem[9][2] ) );
  EDFFX1 \mem_reg[9][1]  ( .D(n883), .E(n981), .CK(clk), .Q(\mem[9][1] ) );
  EDFFX1 \mem_reg[9][0]  ( .D(n877), .E(n981), .CK(clk), .Q(\mem[9][0] ) );
  EDFFX1 \mem_reg[13][7]  ( .D(n919), .E(n990), .CK(clk), .Q(\mem[13][7] ) );
  EDFFX1 \mem_reg[13][6]  ( .D(n913), .E(n990), .CK(clk), .Q(\mem[13][6] ) );
  EDFFX1 \mem_reg[13][5]  ( .D(n907), .E(n990), .CK(clk), .Q(\mem[13][5] ) );
  EDFFX1 \mem_reg[13][4]  ( .D(n901), .E(n990), .CK(clk), .Q(\mem[13][4] ) );
  EDFFX1 \mem_reg[13][3]  ( .D(n895), .E(n990), .CK(clk), .Q(\mem[13][3] ) );
  EDFFX1 \mem_reg[13][2]  ( .D(n889), .E(n990), .CK(clk), .Q(\mem[13][2] ) );
  EDFFX1 \mem_reg[13][1]  ( .D(n883), .E(n990), .CK(clk), .Q(\mem[13][1] ) );
  EDFFX1 \mem_reg[13][0]  ( .D(n877), .E(n990), .CK(clk), .Q(\mem[13][0] ) );
  EDFFX1 \mem_reg[17][7]  ( .D(n919), .E(n962), .CK(clk), .Q(\mem[17][7] ) );
  EDFFX1 \mem_reg[17][6]  ( .D(n913), .E(n962), .CK(clk), .Q(\mem[17][6] ) );
  EDFFX1 \mem_reg[17][5]  ( .D(n907), .E(n962), .CK(clk), .Q(\mem[17][5] ) );
  EDFFX1 \mem_reg[17][4]  ( .D(n901), .E(n962), .CK(clk), .Q(\mem[17][4] ) );
  EDFFX1 \mem_reg[17][3]  ( .D(n895), .E(n962), .CK(clk), .Q(\mem[17][3] ) );
  EDFFX1 \mem_reg[17][2]  ( .D(n889), .E(n962), .CK(clk), .Q(\mem[17][2] ) );
  EDFFX1 \mem_reg[17][1]  ( .D(n883), .E(n962), .CK(clk), .Q(\mem[17][1] ) );
  EDFFX1 \mem_reg[17][0]  ( .D(n877), .E(n962), .CK(clk), .Q(\mem[17][0] ) );
  EDFFX1 \mem_reg[21][7]  ( .D(n918), .E(n971), .CK(clk), .Q(\mem[21][7] ) );
  EDFFX1 \mem_reg[21][6]  ( .D(n912), .E(n971), .CK(clk), .Q(\mem[21][6] ) );
  EDFFX1 \mem_reg[21][5]  ( .D(n906), .E(n971), .CK(clk), .Q(\mem[21][5] ) );
  EDFFX1 \mem_reg[21][4]  ( .D(n900), .E(n971), .CK(clk), .Q(\mem[21][4] ) );
  EDFFX1 \mem_reg[21][3]  ( .D(n894), .E(n971), .CK(clk), .Q(\mem[21][3] ) );
  EDFFX1 \mem_reg[21][2]  ( .D(n888), .E(n971), .CK(clk), .Q(\mem[21][2] ) );
  EDFFX1 \mem_reg[21][1]  ( .D(n882), .E(n971), .CK(clk), .Q(\mem[21][1] ) );
  EDFFX1 \mem_reg[21][0]  ( .D(n876), .E(n971), .CK(clk), .Q(\mem[21][0] ) );
  EDFFX1 \mem_reg[25][7]  ( .D(n918), .E(n980), .CK(clk), .Q(\mem[25][7] ) );
  EDFFX1 \mem_reg[25][6]  ( .D(n912), .E(n980), .CK(clk), .Q(\mem[25][6] ) );
  EDFFX1 \mem_reg[25][5]  ( .D(n906), .E(n980), .CK(clk), .Q(\mem[25][5] ) );
  EDFFX1 \mem_reg[25][4]  ( .D(n900), .E(n980), .CK(clk), .Q(\mem[25][4] ) );
  EDFFX1 \mem_reg[25][3]  ( .D(n894), .E(n980), .CK(clk), .Q(\mem[25][3] ) );
  EDFFX1 \mem_reg[25][2]  ( .D(n888), .E(n980), .CK(clk), .Q(\mem[25][2] ) );
  EDFFX1 \mem_reg[25][1]  ( .D(n882), .E(n980), .CK(clk), .Q(\mem[25][1] ) );
  EDFFX1 \mem_reg[25][0]  ( .D(n876), .E(n980), .CK(clk), .Q(\mem[25][0] ) );
  EDFFX1 \mem_reg[29][7]  ( .D(n918), .E(n989), .CK(clk), .Q(\mem[29][7] ) );
  EDFFX1 \mem_reg[29][6]  ( .D(n912), .E(n989), .CK(clk), .Q(\mem[29][6] ) );
  EDFFX1 \mem_reg[29][5]  ( .D(n906), .E(n989), .CK(clk), .Q(\mem[29][5] ) );
  EDFFX1 \mem_reg[29][4]  ( .D(n900), .E(n989), .CK(clk), .Q(\mem[29][4] ) );
  EDFFX1 \mem_reg[29][3]  ( .D(n894), .E(n989), .CK(clk), .Q(\mem[29][3] ) );
  EDFFX1 \mem_reg[29][2]  ( .D(n888), .E(n989), .CK(clk), .Q(\mem[29][2] ) );
  EDFFX1 \mem_reg[29][1]  ( .D(n882), .E(n989), .CK(clk), .Q(\mem[29][1] ) );
  EDFFX1 \mem_reg[29][0]  ( .D(n876), .E(n989), .CK(clk), .Q(\mem[29][0] ) );
  EDFFX1 \mem_reg[33][7]  ( .D(n917), .E(n961), .CK(clk), .Q(\mem[33][7] ) );
  EDFFX1 \mem_reg[33][6]  ( .D(n911), .E(n961), .CK(clk), .Q(\mem[33][6] ) );
  EDFFX1 \mem_reg[33][5]  ( .D(n905), .E(n961), .CK(clk), .Q(\mem[33][5] ) );
  EDFFX1 \mem_reg[33][4]  ( .D(n899), .E(n961), .CK(clk), .Q(\mem[33][4] ) );
  EDFFX1 \mem_reg[33][3]  ( .D(n893), .E(n961), .CK(clk), .Q(\mem[33][3] ) );
  EDFFX1 \mem_reg[33][2]  ( .D(n887), .E(n961), .CK(clk), .Q(\mem[33][2] ) );
  EDFFX1 \mem_reg[33][1]  ( .D(n881), .E(n961), .CK(clk), .Q(\mem[33][1] ) );
  EDFFX1 \mem_reg[33][0]  ( .D(n875), .E(n961), .CK(clk), .Q(\mem[33][0] ) );
  EDFFX1 \mem_reg[37][7]  ( .D(n917), .E(n970), .CK(clk), .Q(\mem[37][7] ) );
  EDFFX1 \mem_reg[37][6]  ( .D(n911), .E(n970), .CK(clk), .Q(\mem[37][6] ) );
  EDFFX1 \mem_reg[37][5]  ( .D(n905), .E(n970), .CK(clk), .Q(\mem[37][5] ) );
  EDFFX1 \mem_reg[37][4]  ( .D(n899), .E(n970), .CK(clk), .Q(\mem[37][4] ) );
  EDFFX1 \mem_reg[37][3]  ( .D(n893), .E(n970), .CK(clk), .Q(\mem[37][3] ) );
  EDFFX1 \mem_reg[37][2]  ( .D(n887), .E(n970), .CK(clk), .Q(\mem[37][2] ) );
  EDFFX1 \mem_reg[37][1]  ( .D(n881), .E(n970), .CK(clk), .Q(\mem[37][1] ) );
  EDFFX1 \mem_reg[37][0]  ( .D(n875), .E(n970), .CK(clk), .Q(\mem[37][0] ) );
  EDFFX1 \mem_reg[41][7]  ( .D(n917), .E(n979), .CK(clk), .Q(\mem[41][7] ) );
  EDFFX1 \mem_reg[41][6]  ( .D(n911), .E(n979), .CK(clk), .Q(\mem[41][6] ) );
  EDFFX1 \mem_reg[41][5]  ( .D(n905), .E(n979), .CK(clk), .Q(\mem[41][5] ) );
  EDFFX1 \mem_reg[41][4]  ( .D(n899), .E(n979), .CK(clk), .Q(\mem[41][4] ) );
  EDFFX1 \mem_reg[41][3]  ( .D(n893), .E(n979), .CK(clk), .Q(\mem[41][3] ) );
  EDFFX1 \mem_reg[41][2]  ( .D(n887), .E(n979), .CK(clk), .Q(\mem[41][2] ) );
  EDFFX1 \mem_reg[41][1]  ( .D(n881), .E(n979), .CK(clk), .Q(\mem[41][1] ) );
  EDFFX1 \mem_reg[41][0]  ( .D(n875), .E(n979), .CK(clk), .Q(\mem[41][0] ) );
  EDFFX1 \mem_reg[45][7]  ( .D(n916), .E(n988), .CK(clk), .Q(\mem[45][7] ) );
  EDFFX1 \mem_reg[45][6]  ( .D(n910), .E(n988), .CK(clk), .Q(\mem[45][6] ) );
  EDFFX1 \mem_reg[45][5]  ( .D(n904), .E(n988), .CK(clk), .Q(\mem[45][5] ) );
  EDFFX1 \mem_reg[45][4]  ( .D(n898), .E(n988), .CK(clk), .Q(\mem[45][4] ) );
  EDFFX1 \mem_reg[45][3]  ( .D(n892), .E(n988), .CK(clk), .Q(\mem[45][3] ) );
  EDFFX1 \mem_reg[45][2]  ( .D(n886), .E(n988), .CK(clk), .Q(\mem[45][2] ) );
  EDFFX1 \mem_reg[45][1]  ( .D(n880), .E(n988), .CK(clk), .Q(\mem[45][1] ) );
  EDFFX1 \mem_reg[45][0]  ( .D(n874), .E(n988), .CK(clk), .Q(\mem[45][0] ) );
  EDFFX1 \mem_reg[49][7]  ( .D(n916), .E(n960), .CK(clk), .Q(\mem[49][7] ) );
  EDFFX1 \mem_reg[49][6]  ( .D(n910), .E(n960), .CK(clk), .Q(\mem[49][6] ) );
  EDFFX1 \mem_reg[49][5]  ( .D(n904), .E(n960), .CK(clk), .Q(\mem[49][5] ) );
  EDFFX1 \mem_reg[49][4]  ( .D(n898), .E(n960), .CK(clk), .Q(\mem[49][4] ) );
  EDFFX1 \mem_reg[49][3]  ( .D(n892), .E(n960), .CK(clk), .Q(\mem[49][3] ) );
  EDFFX1 \mem_reg[49][2]  ( .D(n886), .E(n960), .CK(clk), .Q(\mem[49][2] ) );
  EDFFX1 \mem_reg[49][1]  ( .D(n880), .E(n960), .CK(clk), .Q(\mem[49][1] ) );
  EDFFX1 \mem_reg[49][0]  ( .D(n874), .E(n960), .CK(clk), .Q(\mem[49][0] ) );
  EDFFX1 \mem_reg[53][7]  ( .D(n916), .E(n969), .CK(clk), .Q(\mem[53][7] ) );
  EDFFX1 \mem_reg[53][6]  ( .D(n910), .E(n969), .CK(clk), .Q(\mem[53][6] ) );
  EDFFX1 \mem_reg[53][5]  ( .D(n904), .E(n969), .CK(clk), .Q(\mem[53][5] ) );
  EDFFX1 \mem_reg[53][4]  ( .D(n898), .E(n969), .CK(clk), .Q(\mem[53][4] ) );
  EDFFX1 \mem_reg[53][3]  ( .D(n892), .E(n969), .CK(clk), .Q(\mem[53][3] ) );
  EDFFX1 \mem_reg[53][2]  ( .D(n886), .E(n969), .CK(clk), .Q(\mem[53][2] ) );
  EDFFX1 \mem_reg[53][1]  ( .D(n880), .E(n969), .CK(clk), .Q(\mem[53][1] ) );
  EDFFX1 \mem_reg[53][0]  ( .D(n874), .E(n969), .CK(clk), .Q(\mem[53][0] ) );
  EDFFX1 \mem_reg[57][7]  ( .D(n915), .E(n978), .CK(clk), .Q(\mem[57][7] ) );
  EDFFX1 \mem_reg[57][6]  ( .D(n909), .E(n978), .CK(clk), .Q(\mem[57][6] ) );
  EDFFX1 \mem_reg[57][5]  ( .D(n903), .E(n978), .CK(clk), .Q(\mem[57][5] ) );
  EDFFX1 \mem_reg[57][4]  ( .D(n897), .E(n978), .CK(clk), .Q(\mem[57][4] ) );
  EDFFX1 \mem_reg[57][3]  ( .D(n891), .E(n978), .CK(clk), .Q(\mem[57][3] ) );
  EDFFX1 \mem_reg[57][2]  ( .D(n885), .E(n978), .CK(clk), .Q(\mem[57][2] ) );
  EDFFX1 \mem_reg[57][1]  ( .D(n879), .E(n978), .CK(clk), .Q(\mem[57][1] ) );
  EDFFX1 \mem_reg[57][0]  ( .D(n873), .E(n978), .CK(clk), .Q(\mem[57][0] ) );
  EDFFX1 \mem_reg[61][7]  ( .D(n918), .E(n987), .CK(clk), .Q(\mem[61][7] ) );
  EDFFX1 \mem_reg[61][6]  ( .D(n912), .E(n987), .CK(clk), .Q(\mem[61][6] ) );
  EDFFX1 \mem_reg[61][5]  ( .D(n906), .E(n987), .CK(clk), .Q(\mem[61][5] ) );
  EDFFX1 \mem_reg[61][4]  ( .D(n900), .E(n987), .CK(clk), .Q(\mem[61][4] ) );
  EDFFX1 \mem_reg[61][3]  ( .D(n894), .E(n987), .CK(clk), .Q(\mem[61][3] ) );
  EDFFX1 \mem_reg[61][2]  ( .D(n888), .E(n987), .CK(clk), .Q(\mem[61][2] ) );
  EDFFX1 \mem_reg[61][1]  ( .D(n882), .E(n987), .CK(clk), .Q(\mem[61][1] ) );
  EDFFX1 \mem_reg[61][0]  ( .D(n876), .E(n987), .CK(clk), .Q(\mem[61][0] ) );
  EDFFX1 \mem_reg[65][7]  ( .D(n916), .E(n959), .CK(clk), .Q(\mem[65][7] ) );
  EDFFX1 \mem_reg[65][6]  ( .D(n910), .E(n959), .CK(clk), .Q(\mem[65][6] ) );
  EDFFX1 \mem_reg[65][5]  ( .D(n904), .E(n959), .CK(clk), .Q(\mem[65][5] ) );
  EDFFX1 \mem_reg[65][4]  ( .D(n898), .E(n959), .CK(clk), .Q(\mem[65][4] ) );
  EDFFX1 \mem_reg[65][3]  ( .D(n892), .E(n959), .CK(clk), .Q(\mem[65][3] ) );
  EDFFX1 \mem_reg[65][2]  ( .D(n886), .E(n959), .CK(clk), .Q(\mem[65][2] ) );
  EDFFX1 \mem_reg[65][1]  ( .D(n880), .E(n959), .CK(clk), .Q(\mem[65][1] ) );
  EDFFX1 \mem_reg[65][0]  ( .D(n874), .E(n959), .CK(clk), .Q(\mem[65][0] ) );
  EDFFX1 \mem_reg[69][7]  ( .D(n915), .E(n968), .CK(clk), .Q(\mem[69][7] ) );
  EDFFX1 \mem_reg[69][6]  ( .D(n909), .E(n968), .CK(clk), .Q(\mem[69][6] ) );
  EDFFX1 \mem_reg[69][5]  ( .D(n903), .E(n968), .CK(clk), .Q(\mem[69][5] ) );
  EDFFX1 \mem_reg[69][4]  ( .D(n897), .E(n968), .CK(clk), .Q(\mem[69][4] ) );
  EDFFX1 \mem_reg[69][3]  ( .D(n891), .E(n968), .CK(clk), .Q(\mem[69][3] ) );
  EDFFX1 \mem_reg[69][2]  ( .D(n885), .E(n968), .CK(clk), .Q(\mem[69][2] ) );
  EDFFX1 \mem_reg[69][1]  ( .D(n879), .E(n968), .CK(clk), .Q(\mem[69][1] ) );
  EDFFX1 \mem_reg[69][0]  ( .D(n873), .E(n968), .CK(clk), .Q(\mem[69][0] ) );
  EDFFX1 \mem_reg[73][7]  ( .D(n915), .E(n977), .CK(clk), .Q(\mem[73][7] ) );
  EDFFX1 \mem_reg[73][6]  ( .D(n909), .E(n977), .CK(clk), .Q(\mem[73][6] ) );
  EDFFX1 \mem_reg[73][5]  ( .D(n903), .E(n977), .CK(clk), .Q(\mem[73][5] ) );
  EDFFX1 \mem_reg[73][4]  ( .D(n897), .E(n977), .CK(clk), .Q(\mem[73][4] ) );
  EDFFX1 \mem_reg[73][3]  ( .D(n891), .E(n977), .CK(clk), .Q(\mem[73][3] ) );
  EDFFX1 \mem_reg[73][2]  ( .D(n885), .E(n977), .CK(clk), .Q(\mem[73][2] ) );
  EDFFX1 \mem_reg[73][1]  ( .D(n879), .E(n977), .CK(clk), .Q(\mem[73][1] ) );
  EDFFX1 \mem_reg[73][0]  ( .D(n873), .E(n977), .CK(clk), .Q(\mem[73][0] ) );
  EDFFX1 \mem_reg[77][7]  ( .D(n915), .E(n986), .CK(clk), .Q(\mem[77][7] ) );
  EDFFX1 \mem_reg[77][6]  ( .D(n909), .E(n986), .CK(clk), .Q(\mem[77][6] ) );
  EDFFX1 \mem_reg[77][5]  ( .D(n903), .E(n986), .CK(clk), .Q(\mem[77][5] ) );
  EDFFX1 \mem_reg[77][4]  ( .D(n897), .E(n986), .CK(clk), .Q(\mem[77][4] ) );
  EDFFX1 \mem_reg[77][3]  ( .D(n891), .E(n986), .CK(clk), .Q(\mem[77][3] ) );
  EDFFX1 \mem_reg[77][2]  ( .D(n885), .E(n986), .CK(clk), .Q(\mem[77][2] ) );
  EDFFX1 \mem_reg[77][1]  ( .D(n879), .E(n986), .CK(clk), .Q(\mem[77][1] ) );
  EDFFX1 \mem_reg[77][0]  ( .D(n873), .E(n986), .CK(clk), .Q(\mem[77][0] ) );
  EDFFX1 \mem_reg[81][7]  ( .D(n914), .E(n958), .CK(clk), .Q(\mem[81][7] ) );
  EDFFX1 \mem_reg[81][6]  ( .D(n908), .E(n958), .CK(clk), .Q(\mem[81][6] ) );
  EDFFX1 \mem_reg[81][5]  ( .D(n902), .E(n958), .CK(clk), .Q(\mem[81][5] ) );
  EDFFX1 \mem_reg[81][4]  ( .D(n896), .E(n958), .CK(clk), .Q(\mem[81][4] ) );
  EDFFX1 \mem_reg[81][3]  ( .D(n890), .E(n958), .CK(clk), .Q(\mem[81][3] ) );
  EDFFX1 \mem_reg[81][2]  ( .D(n884), .E(n958), .CK(clk), .Q(\mem[81][2] ) );
  EDFFX1 \mem_reg[81][1]  ( .D(n878), .E(n958), .CK(clk), .Q(\mem[81][1] ) );
  EDFFX1 \mem_reg[81][0]  ( .D(n872), .E(n958), .CK(clk), .Q(\mem[81][0] ) );
  EDFFX1 \mem_reg[85][7]  ( .D(n914), .E(n967), .CK(clk), .Q(\mem[85][7] ) );
  EDFFX1 \mem_reg[85][6]  ( .D(n908), .E(n967), .CK(clk), .Q(\mem[85][6] ) );
  EDFFX1 \mem_reg[85][5]  ( .D(n902), .E(n967), .CK(clk), .Q(\mem[85][5] ) );
  EDFFX1 \mem_reg[85][4]  ( .D(n896), .E(n967), .CK(clk), .Q(\mem[85][4] ) );
  EDFFX1 \mem_reg[85][3]  ( .D(n890), .E(n967), .CK(clk), .Q(\mem[85][3] ) );
  EDFFX1 \mem_reg[85][2]  ( .D(n884), .E(n967), .CK(clk), .Q(\mem[85][2] ) );
  EDFFX1 \mem_reg[85][1]  ( .D(n878), .E(n967), .CK(clk), .Q(\mem[85][1] ) );
  EDFFX1 \mem_reg[85][0]  ( .D(n872), .E(n967), .CK(clk), .Q(\mem[85][0] ) );
  EDFFX1 \mem_reg[89][7]  ( .D(n914), .E(n976), .CK(clk), .Q(\mem[89][7] ) );
  EDFFX1 \mem_reg[89][6]  ( .D(n908), .E(n976), .CK(clk), .Q(\mem[89][6] ) );
  EDFFX1 \mem_reg[89][5]  ( .D(n902), .E(n976), .CK(clk), .Q(\mem[89][5] ) );
  EDFFX1 \mem_reg[89][4]  ( .D(n896), .E(n976), .CK(clk), .Q(\mem[89][4] ) );
  EDFFX1 \mem_reg[89][3]  ( .D(n890), .E(n976), .CK(clk), .Q(\mem[89][3] ) );
  EDFFX1 \mem_reg[89][2]  ( .D(n884), .E(n976), .CK(clk), .Q(\mem[89][2] ) );
  EDFFX1 \mem_reg[89][1]  ( .D(n878), .E(n976), .CK(clk), .Q(\mem[89][1] ) );
  EDFFX1 \mem_reg[89][0]  ( .D(n872), .E(n976), .CK(clk), .Q(\mem[89][0] ) );
  EDFFX1 \mem_reg[93][7]  ( .D(n915), .E(n985), .CK(clk), .Q(\mem[93][7] ) );
  EDFFX1 \mem_reg[93][6]  ( .D(n909), .E(n985), .CK(clk), .Q(\mem[93][6] ) );
  EDFFX1 \mem_reg[93][5]  ( .D(n903), .E(n985), .CK(clk), .Q(\mem[93][5] ) );
  EDFFX1 \mem_reg[93][4]  ( .D(n897), .E(n985), .CK(clk), .Q(\mem[93][4] ) );
  EDFFX1 \mem_reg[93][3]  ( .D(n891), .E(n985), .CK(clk), .Q(\mem[93][3] ) );
  EDFFX1 \mem_reg[93][2]  ( .D(n885), .E(n985), .CK(clk), .Q(\mem[93][2] ) );
  EDFFX1 \mem_reg[93][1]  ( .D(n879), .E(n985), .CK(clk), .Q(\mem[93][1] ) );
  EDFFX1 \mem_reg[93][0]  ( .D(n873), .E(n985), .CK(clk), .Q(\mem[93][0] ) );
  EDFFX1 \mem_reg[97][7]  ( .D(n914), .E(n957), .CK(clk), .Q(\mem[97][7] ) );
  EDFFX1 \mem_reg[97][6]  ( .D(n908), .E(n957), .CK(clk), .Q(\mem[97][6] ) );
  EDFFX1 \mem_reg[97][5]  ( .D(n902), .E(n957), .CK(clk), .Q(\mem[97][5] ) );
  EDFFX1 \mem_reg[97][4]  ( .D(n896), .E(n957), .CK(clk), .Q(\mem[97][4] ) );
  EDFFX1 \mem_reg[97][3]  ( .D(n890), .E(n957), .CK(clk), .Q(\mem[97][3] ) );
  EDFFX1 \mem_reg[97][2]  ( .D(n884), .E(n957), .CK(clk), .Q(\mem[97][2] ) );
  EDFFX1 \mem_reg[97][1]  ( .D(n878), .E(n957), .CK(clk), .Q(\mem[97][1] ) );
  EDFFX1 \mem_reg[97][0]  ( .D(n872), .E(n957), .CK(clk), .Q(\mem[97][0] ) );
  EDFFX1 \mem_reg[101][7]  ( .D(n915), .E(n966), .CK(clk), .Q(\mem[101][7] )
         );
  EDFFX1 \mem_reg[101][6]  ( .D(n909), .E(n966), .CK(clk), .Q(\mem[101][6] )
         );
  EDFFX1 \mem_reg[101][5]  ( .D(n903), .E(n966), .CK(clk), .Q(\mem[101][5] )
         );
  EDFFX1 \mem_reg[101][4]  ( .D(n897), .E(n966), .CK(clk), .Q(\mem[101][4] )
         );
  EDFFX1 \mem_reg[101][3]  ( .D(n891), .E(n966), .CK(clk), .Q(\mem[101][3] )
         );
  EDFFX1 \mem_reg[101][2]  ( .D(n885), .E(n966), .CK(clk), .Q(\mem[101][2] )
         );
  EDFFX1 \mem_reg[101][1]  ( .D(n879), .E(n966), .CK(clk), .Q(\mem[101][1] )
         );
  EDFFX1 \mem_reg[101][0]  ( .D(n873), .E(n966), .CK(clk), .Q(\mem[101][0] )
         );
  EDFFX1 \mem_reg[105][7]  ( .D(n918), .E(n975), .CK(clk), .Q(\mem[105][7] )
         );
  EDFFX1 \mem_reg[105][6]  ( .D(n912), .E(n975), .CK(clk), .Q(\mem[105][6] )
         );
  EDFFX1 \mem_reg[105][5]  ( .D(n906), .E(n975), .CK(clk), .Q(\mem[105][5] )
         );
  EDFFX1 \mem_reg[105][4]  ( .D(n900), .E(n975), .CK(clk), .Q(\mem[105][4] )
         );
  EDFFX1 \mem_reg[105][3]  ( .D(n894), .E(n975), .CK(clk), .Q(\mem[105][3] )
         );
  EDFFX1 \mem_reg[105][2]  ( .D(n888), .E(n975), .CK(clk), .Q(\mem[105][2] )
         );
  EDFFX1 \mem_reg[105][1]  ( .D(n882), .E(n975), .CK(clk), .Q(\mem[105][1] )
         );
  EDFFX1 \mem_reg[105][0]  ( .D(n876), .E(n975), .CK(clk), .Q(\mem[105][0] )
         );
  EDFFX1 \mem_reg[109][7]  ( .D(n916), .E(n984), .CK(clk), .Q(\mem[109][7] )
         );
  EDFFX1 \mem_reg[109][6]  ( .D(n910), .E(n984), .CK(clk), .Q(\mem[109][6] )
         );
  EDFFX1 \mem_reg[109][5]  ( .D(n904), .E(n984), .CK(clk), .Q(\mem[109][5] )
         );
  EDFFX1 \mem_reg[109][4]  ( .D(n898), .E(n984), .CK(clk), .Q(\mem[109][4] )
         );
  EDFFX1 \mem_reg[109][3]  ( .D(n892), .E(n984), .CK(clk), .Q(\mem[109][3] )
         );
  EDFFX1 \mem_reg[109][2]  ( .D(n886), .E(n984), .CK(clk), .Q(\mem[109][2] )
         );
  EDFFX1 \mem_reg[109][1]  ( .D(n880), .E(n984), .CK(clk), .Q(\mem[109][1] )
         );
  EDFFX1 \mem_reg[109][0]  ( .D(n874), .E(n984), .CK(clk), .Q(\mem[109][0] )
         );
  EDFFX1 \mem_reg[113][7]  ( .D(n919), .E(n956), .CK(clk), .Q(\mem[113][7] )
         );
  EDFFX1 \mem_reg[113][6]  ( .D(n913), .E(n956), .CK(clk), .Q(\mem[113][6] )
         );
  EDFFX1 \mem_reg[113][5]  ( .D(n907), .E(n956), .CK(clk), .Q(\mem[113][5] )
         );
  EDFFX1 \mem_reg[113][4]  ( .D(n901), .E(n956), .CK(clk), .Q(\mem[113][4] )
         );
  EDFFX1 \mem_reg[113][3]  ( .D(n895), .E(n956), .CK(clk), .Q(\mem[113][3] )
         );
  EDFFX1 \mem_reg[113][2]  ( .D(n889), .E(n956), .CK(clk), .Q(\mem[113][2] )
         );
  EDFFX1 \mem_reg[113][1]  ( .D(n883), .E(n956), .CK(clk), .Q(\mem[113][1] )
         );
  EDFFX1 \mem_reg[113][0]  ( .D(n877), .E(n956), .CK(clk), .Q(\mem[113][0] )
         );
  EDFFX1 \mem_reg[117][7]  ( .D(n919), .E(n965), .CK(clk), .Q(\mem[117][7] )
         );
  EDFFX1 \mem_reg[117][6]  ( .D(n913), .E(n965), .CK(clk), .Q(\mem[117][6] )
         );
  EDFFX1 \mem_reg[117][5]  ( .D(n907), .E(n965), .CK(clk), .Q(\mem[117][5] )
         );
  EDFFX1 \mem_reg[117][4]  ( .D(n901), .E(n965), .CK(clk), .Q(\mem[117][4] )
         );
  EDFFX1 \mem_reg[117][3]  ( .D(n895), .E(n965), .CK(clk), .Q(\mem[117][3] )
         );
  EDFFX1 \mem_reg[117][2]  ( .D(n889), .E(n965), .CK(clk), .Q(\mem[117][2] )
         );
  EDFFX1 \mem_reg[117][1]  ( .D(n883), .E(n965), .CK(clk), .Q(\mem[117][1] )
         );
  EDFFX1 \mem_reg[117][0]  ( .D(n877), .E(n965), .CK(clk), .Q(\mem[117][0] )
         );
  EDFFX1 \mem_reg[121][7]  ( .D(n917), .E(n974), .CK(clk), .Q(\mem[121][7] )
         );
  EDFFX1 \mem_reg[121][6]  ( .D(n911), .E(n974), .CK(clk), .Q(\mem[121][6] )
         );
  EDFFX1 \mem_reg[121][5]  ( .D(n905), .E(n974), .CK(clk), .Q(\mem[121][5] )
         );
  EDFFX1 \mem_reg[121][4]  ( .D(n899), .E(n974), .CK(clk), .Q(\mem[121][4] )
         );
  EDFFX1 \mem_reg[121][3]  ( .D(n893), .E(n974), .CK(clk), .Q(\mem[121][3] )
         );
  EDFFX1 \mem_reg[121][2]  ( .D(n887), .E(n974), .CK(clk), .Q(\mem[121][2] )
         );
  EDFFX1 \mem_reg[121][1]  ( .D(n881), .E(n974), .CK(clk), .Q(\mem[121][1] )
         );
  EDFFX1 \mem_reg[121][0]  ( .D(n875), .E(n974), .CK(clk), .Q(\mem[121][0] )
         );
  EDFFX1 \mem_reg[125][7]  ( .D(n918), .E(n983), .CK(clk), .Q(\mem[125][7] )
         );
  EDFFX1 \mem_reg[125][6]  ( .D(n912), .E(n983), .CK(clk), .Q(\mem[125][6] )
         );
  EDFFX1 \mem_reg[125][5]  ( .D(n906), .E(n983), .CK(clk), .Q(\mem[125][5] )
         );
  EDFFX1 \mem_reg[125][4]  ( .D(n900), .E(n983), .CK(clk), .Q(\mem[125][4] )
         );
  EDFFX1 \mem_reg[125][3]  ( .D(n894), .E(n983), .CK(clk), .Q(\mem[125][3] )
         );
  EDFFX1 \mem_reg[125][2]  ( .D(n888), .E(n983), .CK(clk), .Q(\mem[125][2] )
         );
  EDFFX1 \mem_reg[125][1]  ( .D(n882), .E(n983), .CK(clk), .Q(\mem[125][1] )
         );
  EDFFX1 \mem_reg[125][0]  ( .D(n876), .E(n983), .CK(clk), .Q(\mem[125][0] )
         );
  EDFFX1 \mem_reg[3][7]  ( .D(n915), .E(n927), .CK(clk), .Q(\mem[3][7] ) );
  EDFFX1 \mem_reg[3][6]  ( .D(n909), .E(n927), .CK(clk), .Q(\mem[3][6] ) );
  EDFFX1 \mem_reg[3][5]  ( .D(n903), .E(n927), .CK(clk), .Q(\mem[3][5] ) );
  EDFFX1 \mem_reg[3][4]  ( .D(n897), .E(n927), .CK(clk), .Q(\mem[3][4] ) );
  EDFFX1 \mem_reg[3][3]  ( .D(n891), .E(n927), .CK(clk), .Q(\mem[3][3] ) );
  EDFFX1 \mem_reg[3][2]  ( .D(n885), .E(n927), .CK(clk), .Q(\mem[3][2] ) );
  EDFFX1 \mem_reg[3][1]  ( .D(n879), .E(n927), .CK(clk), .Q(\mem[3][1] ) );
  EDFFX1 \mem_reg[3][0]  ( .D(n873), .E(n927), .CK(clk), .Q(\mem[3][0] ) );
  EDFFX1 \mem_reg[7][7]  ( .D(n914), .E(n936), .CK(clk), .Q(\mem[7][7] ) );
  EDFFX1 \mem_reg[7][6]  ( .D(n908), .E(n936), .CK(clk), .Q(\mem[7][6] ) );
  EDFFX1 \mem_reg[7][5]  ( .D(n902), .E(n936), .CK(clk), .Q(\mem[7][5] ) );
  EDFFX1 \mem_reg[7][4]  ( .D(n896), .E(n936), .CK(clk), .Q(\mem[7][4] ) );
  EDFFX1 \mem_reg[7][3]  ( .D(n890), .E(n936), .CK(clk), .Q(\mem[7][3] ) );
  EDFFX1 \mem_reg[7][2]  ( .D(n884), .E(n936), .CK(clk), .Q(\mem[7][2] ) );
  EDFFX1 \mem_reg[7][1]  ( .D(n878), .E(n936), .CK(clk), .Q(\mem[7][1] ) );
  EDFFX1 \mem_reg[7][0]  ( .D(n872), .E(n936), .CK(clk), .Q(\mem[7][0] ) );
  EDFFX1 \mem_reg[11][7]  ( .D(n919), .E(n945), .CK(clk), .Q(\mem[11][7] ) );
  EDFFX1 \mem_reg[11][6]  ( .D(n913), .E(n945), .CK(clk), .Q(\mem[11][6] ) );
  EDFFX1 \mem_reg[11][5]  ( .D(n907), .E(n945), .CK(clk), .Q(\mem[11][5] ) );
  EDFFX1 \mem_reg[11][4]  ( .D(n901), .E(n945), .CK(clk), .Q(\mem[11][4] ) );
  EDFFX1 \mem_reg[11][3]  ( .D(n895), .E(n945), .CK(clk), .Q(\mem[11][3] ) );
  EDFFX1 \mem_reg[11][2]  ( .D(n889), .E(n945), .CK(clk), .Q(\mem[11][2] ) );
  EDFFX1 \mem_reg[11][1]  ( .D(n883), .E(n945), .CK(clk), .Q(\mem[11][1] ) );
  EDFFX1 \mem_reg[11][0]  ( .D(n877), .E(n945), .CK(clk), .Q(\mem[11][0] ) );
  EDFFX1 \mem_reg[15][7]  ( .D(n919), .E(n954), .CK(clk), .Q(\mem[15][7] ) );
  EDFFX1 \mem_reg[15][6]  ( .D(n913), .E(n954), .CK(clk), .Q(\mem[15][6] ) );
  EDFFX1 \mem_reg[15][5]  ( .D(n907), .E(n954), .CK(clk), .Q(\mem[15][5] ) );
  EDFFX1 \mem_reg[15][4]  ( .D(n901), .E(n954), .CK(clk), .Q(\mem[15][4] ) );
  EDFFX1 \mem_reg[15][3]  ( .D(n895), .E(n954), .CK(clk), .Q(\mem[15][3] ) );
  EDFFX1 \mem_reg[15][2]  ( .D(n889), .E(n954), .CK(clk), .Q(\mem[15][2] ) );
  EDFFX1 \mem_reg[15][1]  ( .D(n883), .E(n954), .CK(clk), .Q(\mem[15][1] ) );
  EDFFX1 \mem_reg[15][0]  ( .D(n877), .E(n954), .CK(clk), .Q(\mem[15][0] ) );
  EDFFX1 \mem_reg[19][7]  ( .D(n919), .E(n926), .CK(clk), .Q(\mem[19][7] ) );
  EDFFX1 \mem_reg[19][6]  ( .D(n913), .E(n926), .CK(clk), .Q(\mem[19][6] ) );
  EDFFX1 \mem_reg[19][5]  ( .D(n907), .E(n926), .CK(clk), .Q(\mem[19][5] ) );
  EDFFX1 \mem_reg[19][4]  ( .D(n901), .E(n926), .CK(clk), .Q(\mem[19][4] ) );
  EDFFX1 \mem_reg[19][3]  ( .D(n895), .E(n926), .CK(clk), .Q(\mem[19][3] ) );
  EDFFX1 \mem_reg[19][2]  ( .D(n889), .E(n926), .CK(clk), .Q(\mem[19][2] ) );
  EDFFX1 \mem_reg[19][1]  ( .D(n883), .E(n926), .CK(clk), .Q(\mem[19][1] ) );
  EDFFX1 \mem_reg[19][0]  ( .D(n877), .E(n926), .CK(clk), .Q(\mem[19][0] ) );
  EDFFX1 \mem_reg[23][7]  ( .D(n918), .E(n935), .CK(clk), .Q(\mem[23][7] ) );
  EDFFX1 \mem_reg[23][6]  ( .D(n912), .E(n935), .CK(clk), .Q(\mem[23][6] ) );
  EDFFX1 \mem_reg[23][5]  ( .D(n906), .E(n935), .CK(clk), .Q(\mem[23][5] ) );
  EDFFX1 \mem_reg[23][4]  ( .D(n900), .E(n935), .CK(clk), .Q(\mem[23][4] ) );
  EDFFX1 \mem_reg[23][3]  ( .D(n894), .E(n935), .CK(clk), .Q(\mem[23][3] ) );
  EDFFX1 \mem_reg[23][2]  ( .D(n888), .E(n935), .CK(clk), .Q(\mem[23][2] ) );
  EDFFX1 \mem_reg[23][1]  ( .D(n882), .E(n935), .CK(clk), .Q(\mem[23][1] ) );
  EDFFX1 \mem_reg[23][0]  ( .D(n876), .E(n935), .CK(clk), .Q(\mem[23][0] ) );
  EDFFX1 \mem_reg[27][7]  ( .D(n918), .E(n944), .CK(clk), .Q(\mem[27][7] ) );
  EDFFX1 \mem_reg[27][6]  ( .D(n912), .E(n944), .CK(clk), .Q(\mem[27][6] ) );
  EDFFX1 \mem_reg[27][5]  ( .D(n906), .E(n944), .CK(clk), .Q(\mem[27][5] ) );
  EDFFX1 \mem_reg[27][4]  ( .D(n900), .E(n944), .CK(clk), .Q(\mem[27][4] ) );
  EDFFX1 \mem_reg[27][3]  ( .D(n894), .E(n944), .CK(clk), .Q(\mem[27][3] ) );
  EDFFX1 \mem_reg[27][2]  ( .D(n888), .E(n944), .CK(clk), .Q(\mem[27][2] ) );
  EDFFX1 \mem_reg[27][1]  ( .D(n882), .E(n944), .CK(clk), .Q(\mem[27][1] ) );
  EDFFX1 \mem_reg[27][0]  ( .D(n876), .E(n944), .CK(clk), .Q(\mem[27][0] ) );
  EDFFX1 \mem_reg[31][7]  ( .D(n918), .E(n953), .CK(clk), .Q(\mem[31][7] ) );
  EDFFX1 \mem_reg[31][6]  ( .D(n912), .E(n953), .CK(clk), .Q(\mem[31][6] ) );
  EDFFX1 \mem_reg[31][5]  ( .D(n906), .E(n953), .CK(clk), .Q(\mem[31][5] ) );
  EDFFX1 \mem_reg[31][4]  ( .D(n900), .E(n953), .CK(clk), .Q(\mem[31][4] ) );
  EDFFX1 \mem_reg[31][3]  ( .D(n894), .E(n953), .CK(clk), .Q(\mem[31][3] ) );
  EDFFX1 \mem_reg[31][2]  ( .D(n888), .E(n953), .CK(clk), .Q(\mem[31][2] ) );
  EDFFX1 \mem_reg[31][1]  ( .D(n882), .E(n953), .CK(clk), .Q(\mem[31][1] ) );
  EDFFX1 \mem_reg[31][0]  ( .D(n876), .E(n953), .CK(clk), .Q(\mem[31][0] ) );
  EDFFX1 \mem_reg[35][7]  ( .D(n917), .E(n925), .CK(clk), .Q(\mem[35][7] ) );
  EDFFX1 \mem_reg[35][6]  ( .D(n911), .E(n925), .CK(clk), .Q(\mem[35][6] ) );
  EDFFX1 \mem_reg[35][5]  ( .D(n905), .E(n925), .CK(clk), .Q(\mem[35][5] ) );
  EDFFX1 \mem_reg[35][4]  ( .D(n899), .E(n925), .CK(clk), .Q(\mem[35][4] ) );
  EDFFX1 \mem_reg[35][3]  ( .D(n893), .E(n925), .CK(clk), .Q(\mem[35][3] ) );
  EDFFX1 \mem_reg[35][2]  ( .D(n887), .E(n925), .CK(clk), .Q(\mem[35][2] ) );
  EDFFX1 \mem_reg[35][1]  ( .D(n881), .E(n925), .CK(clk), .Q(\mem[35][1] ) );
  EDFFX1 \mem_reg[35][0]  ( .D(n875), .E(n925), .CK(clk), .Q(\mem[35][0] ) );
  EDFFX1 \mem_reg[39][7]  ( .D(n917), .E(n934), .CK(clk), .Q(\mem[39][7] ) );
  EDFFX1 \mem_reg[39][6]  ( .D(n911), .E(n934), .CK(clk), .Q(\mem[39][6] ) );
  EDFFX1 \mem_reg[39][5]  ( .D(n905), .E(n934), .CK(clk), .Q(\mem[39][5] ) );
  EDFFX1 \mem_reg[39][4]  ( .D(n899), .E(n934), .CK(clk), .Q(\mem[39][4] ) );
  EDFFX1 \mem_reg[39][3]  ( .D(n893), .E(n934), .CK(clk), .Q(\mem[39][3] ) );
  EDFFX1 \mem_reg[39][2]  ( .D(n887), .E(n934), .CK(clk), .Q(\mem[39][2] ) );
  EDFFX1 \mem_reg[39][1]  ( .D(n881), .E(n934), .CK(clk), .Q(\mem[39][1] ) );
  EDFFX1 \mem_reg[39][0]  ( .D(n875), .E(n934), .CK(clk), .Q(\mem[39][0] ) );
  EDFFX1 \mem_reg[43][7]  ( .D(n917), .E(n943), .CK(clk), .Q(\mem[43][7] ) );
  EDFFX1 \mem_reg[43][6]  ( .D(n911), .E(n943), .CK(clk), .Q(\mem[43][6] ) );
  EDFFX1 \mem_reg[43][5]  ( .D(n905), .E(n943), .CK(clk), .Q(\mem[43][5] ) );
  EDFFX1 \mem_reg[43][4]  ( .D(n899), .E(n943), .CK(clk), .Q(\mem[43][4] ) );
  EDFFX1 \mem_reg[43][3]  ( .D(n893), .E(n943), .CK(clk), .Q(\mem[43][3] ) );
  EDFFX1 \mem_reg[43][2]  ( .D(n887), .E(n943), .CK(clk), .Q(\mem[43][2] ) );
  EDFFX1 \mem_reg[43][1]  ( .D(n881), .E(n943), .CK(clk), .Q(\mem[43][1] ) );
  EDFFX1 \mem_reg[43][0]  ( .D(n875), .E(n943), .CK(clk), .Q(\mem[43][0] ) );
  EDFFX1 \mem_reg[47][7]  ( .D(n916), .E(n952), .CK(clk), .Q(\mem[47][7] ) );
  EDFFX1 \mem_reg[47][6]  ( .D(n910), .E(n952), .CK(clk), .Q(\mem[47][6] ) );
  EDFFX1 \mem_reg[47][5]  ( .D(n904), .E(n952), .CK(clk), .Q(\mem[47][5] ) );
  EDFFX1 \mem_reg[47][4]  ( .D(n898), .E(n952), .CK(clk), .Q(\mem[47][4] ) );
  EDFFX1 \mem_reg[47][3]  ( .D(n892), .E(n952), .CK(clk), .Q(\mem[47][3] ) );
  EDFFX1 \mem_reg[47][2]  ( .D(n886), .E(n952), .CK(clk), .Q(\mem[47][2] ) );
  EDFFX1 \mem_reg[47][1]  ( .D(n880), .E(n952), .CK(clk), .Q(\mem[47][1] ) );
  EDFFX1 \mem_reg[47][0]  ( .D(n874), .E(n952), .CK(clk), .Q(\mem[47][0] ) );
  EDFFX1 \mem_reg[51][7]  ( .D(n916), .E(n924), .CK(clk), .Q(\mem[51][7] ) );
  EDFFX1 \mem_reg[51][6]  ( .D(n910), .E(n924), .CK(clk), .Q(\mem[51][6] ) );
  EDFFX1 \mem_reg[51][5]  ( .D(n904), .E(n924), .CK(clk), .Q(\mem[51][5] ) );
  EDFFX1 \mem_reg[51][4]  ( .D(n898), .E(n924), .CK(clk), .Q(\mem[51][4] ) );
  EDFFX1 \mem_reg[51][3]  ( .D(n892), .E(n924), .CK(clk), .Q(\mem[51][3] ) );
  EDFFX1 \mem_reg[51][2]  ( .D(n886), .E(n924), .CK(clk), .Q(\mem[51][2] ) );
  EDFFX1 \mem_reg[51][1]  ( .D(n880), .E(n924), .CK(clk), .Q(\mem[51][1] ) );
  EDFFX1 \mem_reg[51][0]  ( .D(n874), .E(n924), .CK(clk), .Q(\mem[51][0] ) );
  EDFFX1 \mem_reg[55][7]  ( .D(n916), .E(n933), .CK(clk), .Q(\mem[55][7] ) );
  EDFFX1 \mem_reg[55][6]  ( .D(n910), .E(n933), .CK(clk), .Q(\mem[55][6] ) );
  EDFFX1 \mem_reg[55][5]  ( .D(n904), .E(n933), .CK(clk), .Q(\mem[55][5] ) );
  EDFFX1 \mem_reg[55][4]  ( .D(n898), .E(n933), .CK(clk), .Q(\mem[55][4] ) );
  EDFFX1 \mem_reg[55][3]  ( .D(n892), .E(n933), .CK(clk), .Q(\mem[55][3] ) );
  EDFFX1 \mem_reg[55][2]  ( .D(n886), .E(n933), .CK(clk), .Q(\mem[55][2] ) );
  EDFFX1 \mem_reg[55][1]  ( .D(n880), .E(n933), .CK(clk), .Q(\mem[55][1] ) );
  EDFFX1 \mem_reg[55][0]  ( .D(n874), .E(n933), .CK(clk), .Q(\mem[55][0] ) );
  EDFFX1 \mem_reg[59][7]  ( .D(n919), .E(n942), .CK(clk), .Q(\mem[59][7] ) );
  EDFFX1 \mem_reg[59][6]  ( .D(n913), .E(n942), .CK(clk), .Q(\mem[59][6] ) );
  EDFFX1 \mem_reg[59][5]  ( .D(n907), .E(n942), .CK(clk), .Q(\mem[59][5] ) );
  EDFFX1 \mem_reg[59][4]  ( .D(n901), .E(n942), .CK(clk), .Q(\mem[59][4] ) );
  EDFFX1 \mem_reg[59][3]  ( .D(n895), .E(n942), .CK(clk), .Q(\mem[59][3] ) );
  EDFFX1 \mem_reg[59][2]  ( .D(n889), .E(n942), .CK(clk), .Q(\mem[59][2] ) );
  EDFFX1 \mem_reg[59][1]  ( .D(n883), .E(n942), .CK(clk), .Q(\mem[59][1] ) );
  EDFFX1 \mem_reg[59][0]  ( .D(n877), .E(n942), .CK(clk), .Q(\mem[59][0] ) );
  EDFFX1 \mem_reg[63][7]  ( .D(n917), .E(n951), .CK(clk), .Q(\mem[63][7] ) );
  EDFFX1 \mem_reg[63][6]  ( .D(n911), .E(n951), .CK(clk), .Q(\mem[63][6] ) );
  EDFFX1 \mem_reg[63][5]  ( .D(n905), .E(n951), .CK(clk), .Q(\mem[63][5] ) );
  EDFFX1 \mem_reg[63][4]  ( .D(n899), .E(n951), .CK(clk), .Q(\mem[63][4] ) );
  EDFFX1 \mem_reg[63][3]  ( .D(n893), .E(n951), .CK(clk), .Q(\mem[63][3] ) );
  EDFFX1 \mem_reg[63][2]  ( .D(n887), .E(n951), .CK(clk), .Q(\mem[63][2] ) );
  EDFFX1 \mem_reg[63][1]  ( .D(n881), .E(n951), .CK(clk), .Q(\mem[63][1] ) );
  EDFFX1 \mem_reg[63][0]  ( .D(n875), .E(n951), .CK(clk), .Q(\mem[63][0] ) );
  EDFFX1 \mem_reg[67][7]  ( .D(n916), .E(n923), .CK(clk), .Q(\mem[67][7] ) );
  EDFFX1 \mem_reg[67][6]  ( .D(n910), .E(n923), .CK(clk), .Q(\mem[67][6] ) );
  EDFFX1 \mem_reg[67][5]  ( .D(n904), .E(n923), .CK(clk), .Q(\mem[67][5] ) );
  EDFFX1 \mem_reg[67][4]  ( .D(n898), .E(n923), .CK(clk), .Q(\mem[67][4] ) );
  EDFFX1 \mem_reg[67][3]  ( .D(n892), .E(n923), .CK(clk), .Q(\mem[67][3] ) );
  EDFFX1 \mem_reg[67][2]  ( .D(n886), .E(n923), .CK(clk), .Q(\mem[67][2] ) );
  EDFFX1 \mem_reg[67][1]  ( .D(n880), .E(n923), .CK(clk), .Q(\mem[67][1] ) );
  EDFFX1 \mem_reg[67][0]  ( .D(n874), .E(n923), .CK(clk), .Q(\mem[67][0] ) );
  EDFFX1 \mem_reg[71][7]  ( .D(n915), .E(n932), .CK(clk), .Q(\mem[71][7] ) );
  EDFFX1 \mem_reg[71][6]  ( .D(n909), .E(n932), .CK(clk), .Q(\mem[71][6] ) );
  EDFFX1 \mem_reg[71][5]  ( .D(n903), .E(n932), .CK(clk), .Q(\mem[71][5] ) );
  EDFFX1 \mem_reg[71][4]  ( .D(n897), .E(n932), .CK(clk), .Q(\mem[71][4] ) );
  EDFFX1 \mem_reg[71][3]  ( .D(n891), .E(n932), .CK(clk), .Q(\mem[71][3] ) );
  EDFFX1 \mem_reg[71][2]  ( .D(n885), .E(n932), .CK(clk), .Q(\mem[71][2] ) );
  EDFFX1 \mem_reg[71][1]  ( .D(n879), .E(n932), .CK(clk), .Q(\mem[71][1] ) );
  EDFFX1 \mem_reg[71][0]  ( .D(n873), .E(n932), .CK(clk), .Q(\mem[71][0] ) );
  EDFFX1 \mem_reg[75][7]  ( .D(n915), .E(n941), .CK(clk), .Q(\mem[75][7] ) );
  EDFFX1 \mem_reg[75][6]  ( .D(n909), .E(n941), .CK(clk), .Q(\mem[75][6] ) );
  EDFFX1 \mem_reg[75][5]  ( .D(n903), .E(n941), .CK(clk), .Q(\mem[75][5] ) );
  EDFFX1 \mem_reg[75][4]  ( .D(n897), .E(n941), .CK(clk), .Q(\mem[75][4] ) );
  EDFFX1 \mem_reg[75][3]  ( .D(n891), .E(n941), .CK(clk), .Q(\mem[75][3] ) );
  EDFFX1 \mem_reg[75][2]  ( .D(n885), .E(n941), .CK(clk), .Q(\mem[75][2] ) );
  EDFFX1 \mem_reg[75][1]  ( .D(n879), .E(n941), .CK(clk), .Q(\mem[75][1] ) );
  EDFFX1 \mem_reg[75][0]  ( .D(n873), .E(n941), .CK(clk), .Q(\mem[75][0] ) );
  EDFFX1 \mem_reg[79][7]  ( .D(n915), .E(n950), .CK(clk), .Q(\mem[79][7] ) );
  EDFFX1 \mem_reg[79][6]  ( .D(n909), .E(n950), .CK(clk), .Q(\mem[79][6] ) );
  EDFFX1 \mem_reg[79][5]  ( .D(n903), .E(n950), .CK(clk), .Q(\mem[79][5] ) );
  EDFFX1 \mem_reg[79][4]  ( .D(n897), .E(n950), .CK(clk), .Q(\mem[79][4] ) );
  EDFFX1 \mem_reg[79][3]  ( .D(n891), .E(n950), .CK(clk), .Q(\mem[79][3] ) );
  EDFFX1 \mem_reg[79][2]  ( .D(n885), .E(n950), .CK(clk), .Q(\mem[79][2] ) );
  EDFFX1 \mem_reg[79][1]  ( .D(n879), .E(n950), .CK(clk), .Q(\mem[79][1] ) );
  EDFFX1 \mem_reg[79][0]  ( .D(n873), .E(n950), .CK(clk), .Q(\mem[79][0] ) );
  EDFFX1 \mem_reg[83][7]  ( .D(n914), .E(n922), .CK(clk), .Q(\mem[83][7] ) );
  EDFFX1 \mem_reg[83][6]  ( .D(n908), .E(n922), .CK(clk), .Q(\mem[83][6] ) );
  EDFFX1 \mem_reg[83][5]  ( .D(n902), .E(n922), .CK(clk), .Q(\mem[83][5] ) );
  EDFFX1 \mem_reg[83][4]  ( .D(n896), .E(n922), .CK(clk), .Q(\mem[83][4] ) );
  EDFFX1 \mem_reg[83][3]  ( .D(n890), .E(n922), .CK(clk), .Q(\mem[83][3] ) );
  EDFFX1 \mem_reg[83][2]  ( .D(n884), .E(n922), .CK(clk), .Q(\mem[83][2] ) );
  EDFFX1 \mem_reg[83][1]  ( .D(n878), .E(n922), .CK(clk), .Q(\mem[83][1] ) );
  EDFFX1 \mem_reg[83][0]  ( .D(n872), .E(n922), .CK(clk), .Q(\mem[83][0] ) );
  EDFFX1 \mem_reg[87][7]  ( .D(n914), .E(n931), .CK(clk), .Q(\mem[87][7] ) );
  EDFFX1 \mem_reg[87][6]  ( .D(n908), .E(n931), .CK(clk), .Q(\mem[87][6] ) );
  EDFFX1 \mem_reg[87][5]  ( .D(n902), .E(n931), .CK(clk), .Q(\mem[87][5] ) );
  EDFFX1 \mem_reg[87][4]  ( .D(n896), .E(n931), .CK(clk), .Q(\mem[87][4] ) );
  EDFFX1 \mem_reg[87][3]  ( .D(n890), .E(n931), .CK(clk), .Q(\mem[87][3] ) );
  EDFFX1 \mem_reg[87][2]  ( .D(n884), .E(n931), .CK(clk), .Q(\mem[87][2] ) );
  EDFFX1 \mem_reg[87][1]  ( .D(n878), .E(n931), .CK(clk), .Q(\mem[87][1] ) );
  EDFFX1 \mem_reg[87][0]  ( .D(n872), .E(n931), .CK(clk), .Q(\mem[87][0] ) );
  EDFFX1 \mem_reg[91][7]  ( .D(n914), .E(n940), .CK(clk), .Q(\mem[91][7] ) );
  EDFFX1 \mem_reg[91][6]  ( .D(n908), .E(n940), .CK(clk), .Q(\mem[91][6] ) );
  EDFFX1 \mem_reg[91][5]  ( .D(n902), .E(n940), .CK(clk), .Q(\mem[91][5] ) );
  EDFFX1 \mem_reg[91][4]  ( .D(n896), .E(n940), .CK(clk), .Q(\mem[91][4] ) );
  EDFFX1 \mem_reg[91][3]  ( .D(n890), .E(n940), .CK(clk), .Q(\mem[91][3] ) );
  EDFFX1 \mem_reg[91][2]  ( .D(n884), .E(n940), .CK(clk), .Q(\mem[91][2] ) );
  EDFFX1 \mem_reg[91][1]  ( .D(n878), .E(n940), .CK(clk), .Q(\mem[91][1] ) );
  EDFFX1 \mem_reg[91][0]  ( .D(n872), .E(n940), .CK(clk), .Q(\mem[91][0] ) );
  EDFFX1 \mem_reg[95][7]  ( .D(n919), .E(n949), .CK(clk), .Q(\mem[95][7] ) );
  EDFFX1 \mem_reg[95][6]  ( .D(n913), .E(n949), .CK(clk), .Q(\mem[95][6] ) );
  EDFFX1 \mem_reg[95][5]  ( .D(n907), .E(n949), .CK(clk), .Q(\mem[95][5] ) );
  EDFFX1 \mem_reg[95][4]  ( .D(n901), .E(n949), .CK(clk), .Q(\mem[95][4] ) );
  EDFFX1 \mem_reg[95][3]  ( .D(n895), .E(n949), .CK(clk), .Q(\mem[95][3] ) );
  EDFFX1 \mem_reg[95][2]  ( .D(n889), .E(n949), .CK(clk), .Q(\mem[95][2] ) );
  EDFFX1 \mem_reg[95][1]  ( .D(n883), .E(n949), .CK(clk), .Q(\mem[95][1] ) );
  EDFFX1 \mem_reg[95][0]  ( .D(n877), .E(n949), .CK(clk), .Q(\mem[95][0] ) );
  EDFFX1 \mem_reg[99][7]  ( .D(n914), .E(n921), .CK(clk), .Q(\mem[99][7] ) );
  EDFFX1 \mem_reg[99][6]  ( .D(n908), .E(n921), .CK(clk), .Q(\mem[99][6] ) );
  EDFFX1 \mem_reg[99][5]  ( .D(n902), .E(n921), .CK(clk), .Q(\mem[99][5] ) );
  EDFFX1 \mem_reg[99][4]  ( .D(n896), .E(n921), .CK(clk), .Q(\mem[99][4] ) );
  EDFFX1 \mem_reg[99][3]  ( .D(n890), .E(n921), .CK(clk), .Q(\mem[99][3] ) );
  EDFFX1 \mem_reg[99][2]  ( .D(n884), .E(n921), .CK(clk), .Q(\mem[99][2] ) );
  EDFFX1 \mem_reg[99][1]  ( .D(n878), .E(n921), .CK(clk), .Q(\mem[99][1] ) );
  EDFFX1 \mem_reg[99][0]  ( .D(n872), .E(n921), .CK(clk), .Q(\mem[99][0] ) );
  EDFFX1 \mem_reg[103][7]  ( .D(n917), .E(n930), .CK(clk), .Q(\mem[103][7] )
         );
  EDFFX1 \mem_reg[103][6]  ( .D(n911), .E(n930), .CK(clk), .Q(\mem[103][6] )
         );
  EDFFX1 \mem_reg[103][5]  ( .D(n905), .E(n930), .CK(clk), .Q(\mem[103][5] )
         );
  EDFFX1 \mem_reg[103][4]  ( .D(n899), .E(n930), .CK(clk), .Q(\mem[103][4] )
         );
  EDFFX1 \mem_reg[103][3]  ( .D(n893), .E(n930), .CK(clk), .Q(\mem[103][3] )
         );
  EDFFX1 \mem_reg[103][2]  ( .D(n887), .E(n930), .CK(clk), .Q(\mem[103][2] )
         );
  EDFFX1 \mem_reg[103][1]  ( .D(n881), .E(n930), .CK(clk), .Q(\mem[103][1] )
         );
  EDFFX1 \mem_reg[103][0]  ( .D(n875), .E(n930), .CK(clk), .Q(\mem[103][0] )
         );
  EDFFX1 \mem_reg[107][7]  ( .D(n919), .E(n939), .CK(clk), .Q(\mem[107][7] )
         );
  EDFFX1 \mem_reg[107][6]  ( .D(n913), .E(n939), .CK(clk), .Q(\mem[107][6] )
         );
  EDFFX1 \mem_reg[107][5]  ( .D(n907), .E(n939), .CK(clk), .Q(\mem[107][5] )
         );
  EDFFX1 \mem_reg[107][4]  ( .D(n901), .E(n939), .CK(clk), .Q(\mem[107][4] )
         );
  EDFFX1 \mem_reg[107][3]  ( .D(n895), .E(n939), .CK(clk), .Q(\mem[107][3] )
         );
  EDFFX1 \mem_reg[107][2]  ( .D(n889), .E(n939), .CK(clk), .Q(\mem[107][2] )
         );
  EDFFX1 \mem_reg[107][1]  ( .D(n883), .E(n939), .CK(clk), .Q(\mem[107][1] )
         );
  EDFFX1 \mem_reg[107][0]  ( .D(n877), .E(n939), .CK(clk), .Q(\mem[107][0] )
         );
  EDFFX1 \mem_reg[111][7]  ( .D(n917), .E(n948), .CK(clk), .Q(\mem[111][7] )
         );
  EDFFX1 \mem_reg[111][6]  ( .D(n911), .E(n948), .CK(clk), .Q(\mem[111][6] )
         );
  EDFFX1 \mem_reg[111][5]  ( .D(n905), .E(n948), .CK(clk), .Q(\mem[111][5] )
         );
  EDFFX1 \mem_reg[111][4]  ( .D(n899), .E(n948), .CK(clk), .Q(\mem[111][4] )
         );
  EDFFX1 \mem_reg[111][3]  ( .D(n893), .E(n948), .CK(clk), .Q(\mem[111][3] )
         );
  EDFFX1 \mem_reg[111][2]  ( .D(n887), .E(n948), .CK(clk), .Q(\mem[111][2] )
         );
  EDFFX1 \mem_reg[111][1]  ( .D(n881), .E(n948), .CK(clk), .Q(\mem[111][1] )
         );
  EDFFX1 \mem_reg[111][0]  ( .D(n875), .E(n948), .CK(clk), .Q(\mem[111][0] )
         );
  EDFFX1 \mem_reg[115][7]  ( .D(n918), .E(n920), .CK(clk), .Q(\mem[115][7] )
         );
  EDFFX1 \mem_reg[115][6]  ( .D(n912), .E(n920), .CK(clk), .Q(\mem[115][6] )
         );
  EDFFX1 \mem_reg[115][5]  ( .D(n906), .E(n920), .CK(clk), .Q(\mem[115][5] )
         );
  EDFFX1 \mem_reg[115][4]  ( .D(n900), .E(n920), .CK(clk), .Q(\mem[115][4] )
         );
  EDFFX1 \mem_reg[115][3]  ( .D(n894), .E(n920), .CK(clk), .Q(\mem[115][3] )
         );
  EDFFX1 \mem_reg[115][2]  ( .D(n888), .E(n920), .CK(clk), .Q(\mem[115][2] )
         );
  EDFFX1 \mem_reg[115][1]  ( .D(n882), .E(n920), .CK(clk), .Q(\mem[115][1] )
         );
  EDFFX1 \mem_reg[115][0]  ( .D(n876), .E(n920), .CK(clk), .Q(\mem[115][0] )
         );
  EDFFX1 \mem_reg[119][7]  ( .D(n916), .E(n929), .CK(clk), .Q(\mem[119][7] )
         );
  EDFFX1 \mem_reg[119][6]  ( .D(n910), .E(n929), .CK(clk), .Q(\mem[119][6] )
         );
  EDFFX1 \mem_reg[119][5]  ( .D(n904), .E(n929), .CK(clk), .Q(\mem[119][5] )
         );
  EDFFX1 \mem_reg[119][4]  ( .D(n898), .E(n929), .CK(clk), .Q(\mem[119][4] )
         );
  EDFFX1 \mem_reg[119][3]  ( .D(n892), .E(n929), .CK(clk), .Q(\mem[119][3] )
         );
  EDFFX1 \mem_reg[119][2]  ( .D(n886), .E(n929), .CK(clk), .Q(\mem[119][2] )
         );
  EDFFX1 \mem_reg[119][1]  ( .D(n880), .E(n929), .CK(clk), .Q(\mem[119][1] )
         );
  EDFFX1 \mem_reg[119][0]  ( .D(n874), .E(n929), .CK(clk), .Q(\mem[119][0] )
         );
  EDFFX1 \mem_reg[123][7]  ( .D(n919), .E(n938), .CK(clk), .Q(\mem[123][7] )
         );
  EDFFX1 \mem_reg[123][6]  ( .D(n913), .E(n938), .CK(clk), .Q(\mem[123][6] )
         );
  EDFFX1 \mem_reg[123][5]  ( .D(n907), .E(n938), .CK(clk), .Q(\mem[123][5] )
         );
  EDFFX1 \mem_reg[123][4]  ( .D(n901), .E(n938), .CK(clk), .Q(\mem[123][4] )
         );
  EDFFX1 \mem_reg[123][3]  ( .D(n895), .E(n938), .CK(clk), .Q(\mem[123][3] )
         );
  EDFFX1 \mem_reg[123][2]  ( .D(n889), .E(n938), .CK(clk), .Q(\mem[123][2] )
         );
  EDFFX1 \mem_reg[123][1]  ( .D(n883), .E(n938), .CK(clk), .Q(\mem[123][1] )
         );
  EDFFX1 \mem_reg[123][0]  ( .D(n877), .E(n938), .CK(clk), .Q(\mem[123][0] )
         );
  EDFFX1 \mem_reg[127][7]  ( .D(n917), .E(n947), .CK(clk), .Q(\mem[127][7] )
         );
  EDFFX1 \mem_reg[127][6]  ( .D(n911), .E(n947), .CK(clk), .Q(\mem[127][6] )
         );
  EDFFX1 \mem_reg[127][5]  ( .D(n905), .E(n947), .CK(clk), .Q(\mem[127][5] )
         );
  EDFFX1 \mem_reg[127][4]  ( .D(n899), .E(n947), .CK(clk), .Q(\mem[127][4] )
         );
  EDFFX1 \mem_reg[127][3]  ( .D(n893), .E(n947), .CK(clk), .Q(\mem[127][3] )
         );
  EDFFX1 \mem_reg[127][2]  ( .D(n887), .E(n947), .CK(clk), .Q(\mem[127][2] )
         );
  EDFFX1 \mem_reg[127][1]  ( .D(n881), .E(n947), .CK(clk), .Q(\mem[127][1] )
         );
  EDFFX1 \mem_reg[127][0]  ( .D(n875), .E(n947), .CK(clk), .Q(\mem[127][0] )
         );
  EDFFX1 \mem_reg[0][7]  ( .D(n915), .E(n1000), .CK(clk), .Q(\mem[0][7] ) );
  EDFFX1 \mem_reg[0][6]  ( .D(n909), .E(n1000), .CK(clk), .Q(\mem[0][6] ) );
  EDFFX1 \mem_reg[0][5]  ( .D(n903), .E(n1000), .CK(clk), .Q(\mem[0][5] ) );
  EDFFX1 \mem_reg[0][4]  ( .D(n897), .E(n1000), .CK(clk), .Q(\mem[0][4] ) );
  EDFFX1 \mem_reg[0][3]  ( .D(n891), .E(n1000), .CK(clk), .Q(\mem[0][3] ) );
  EDFFX1 \mem_reg[0][2]  ( .D(n885), .E(n1000), .CK(clk), .Q(\mem[0][2] ) );
  EDFFX1 \mem_reg[0][1]  ( .D(n879), .E(n1000), .CK(clk), .Q(\mem[0][1] ) );
  EDFFX1 \mem_reg[0][0]  ( .D(n873), .E(n1000), .CK(clk), .Q(\mem[0][0] ) );
  EDFFX1 \mem_reg[4][7]  ( .D(n914), .E(n1009), .CK(clk), .Q(\mem[4][7] ) );
  EDFFX1 \mem_reg[4][6]  ( .D(n908), .E(n1009), .CK(clk), .Q(\mem[4][6] ) );
  EDFFX1 \mem_reg[4][5]  ( .D(n902), .E(n1009), .CK(clk), .Q(\mem[4][5] ) );
  EDFFX1 \mem_reg[4][4]  ( .D(n896), .E(n1009), .CK(clk), .Q(\mem[4][4] ) );
  EDFFX1 \mem_reg[4][3]  ( .D(n890), .E(n1009), .CK(clk), .Q(\mem[4][3] ) );
  EDFFX1 \mem_reg[4][2]  ( .D(n884), .E(n1009), .CK(clk), .Q(\mem[4][2] ) );
  EDFFX1 \mem_reg[4][1]  ( .D(n878), .E(n1009), .CK(clk), .Q(\mem[4][1] ) );
  EDFFX1 \mem_reg[4][0]  ( .D(n872), .E(n1009), .CK(clk), .Q(\mem[4][0] ) );
  EDFFX1 \mem_reg[8][7]  ( .D(n919), .E(n1018), .CK(clk), .Q(\mem[8][7] ) );
  EDFFX1 \mem_reg[8][6]  ( .D(n913), .E(n1018), .CK(clk), .Q(\mem[8][6] ) );
  EDFFX1 \mem_reg[8][5]  ( .D(n907), .E(n1018), .CK(clk), .Q(\mem[8][5] ) );
  EDFFX1 \mem_reg[8][4]  ( .D(n901), .E(n1018), .CK(clk), .Q(\mem[8][4] ) );
  EDFFX1 \mem_reg[8][3]  ( .D(n895), .E(n1018), .CK(clk), .Q(\mem[8][3] ) );
  EDFFX1 \mem_reg[8][2]  ( .D(n889), .E(n1018), .CK(clk), .Q(\mem[8][2] ) );
  EDFFX1 \mem_reg[8][1]  ( .D(n883), .E(n1018), .CK(clk), .Q(\mem[8][1] ) );
  EDFFX1 \mem_reg[8][0]  ( .D(n877), .E(n1018), .CK(clk), .Q(\mem[8][0] ) );
  EDFFX1 \mem_reg[12][7]  ( .D(n919), .E(n1027), .CK(clk), .Q(\mem[12][7] ) );
  EDFFX1 \mem_reg[12][6]  ( .D(n913), .E(n1027), .CK(clk), .Q(\mem[12][6] ) );
  EDFFX1 \mem_reg[12][5]  ( .D(n907), .E(n1027), .CK(clk), .Q(\mem[12][5] ) );
  EDFFX1 \mem_reg[12][4]  ( .D(n901), .E(n1027), .CK(clk), .Q(\mem[12][4] ) );
  EDFFX1 \mem_reg[12][3]  ( .D(n895), .E(n1027), .CK(clk), .Q(\mem[12][3] ) );
  EDFFX1 \mem_reg[12][2]  ( .D(n889), .E(n1027), .CK(clk), .Q(\mem[12][2] ) );
  EDFFX1 \mem_reg[12][1]  ( .D(n883), .E(n1027), .CK(clk), .Q(\mem[12][1] ) );
  EDFFX1 \mem_reg[12][0]  ( .D(n877), .E(n1027), .CK(clk), .Q(\mem[12][0] ) );
  EDFFX1 \mem_reg[16][7]  ( .D(n919), .E(n999), .CK(clk), .Q(\mem[16][7] ) );
  EDFFX1 \mem_reg[16][6]  ( .D(n913), .E(n999), .CK(clk), .Q(\mem[16][6] ) );
  EDFFX1 \mem_reg[16][5]  ( .D(n907), .E(n999), .CK(clk), .Q(\mem[16][5] ) );
  EDFFX1 \mem_reg[16][4]  ( .D(n901), .E(n999), .CK(clk), .Q(\mem[16][4] ) );
  EDFFX1 \mem_reg[16][3]  ( .D(n895), .E(n999), .CK(clk), .Q(\mem[16][3] ) );
  EDFFX1 \mem_reg[16][2]  ( .D(n889), .E(n999), .CK(clk), .Q(\mem[16][2] ) );
  EDFFX1 \mem_reg[16][1]  ( .D(n883), .E(n999), .CK(clk), .Q(\mem[16][1] ) );
  EDFFX1 \mem_reg[16][0]  ( .D(n877), .E(n999), .CK(clk), .Q(\mem[16][0] ) );
  EDFFX1 \mem_reg[20][7]  ( .D(n918), .E(n1008), .CK(clk), .Q(\mem[20][7] ) );
  EDFFX1 \mem_reg[20][6]  ( .D(n912), .E(n1008), .CK(clk), .Q(\mem[20][6] ) );
  EDFFX1 \mem_reg[20][5]  ( .D(n906), .E(n1008), .CK(clk), .Q(\mem[20][5] ) );
  EDFFX1 \mem_reg[20][4]  ( .D(n900), .E(n1008), .CK(clk), .Q(\mem[20][4] ) );
  EDFFX1 \mem_reg[20][3]  ( .D(n894), .E(n1008), .CK(clk), .Q(\mem[20][3] ) );
  EDFFX1 \mem_reg[20][2]  ( .D(n888), .E(n1008), .CK(clk), .Q(\mem[20][2] ) );
  EDFFX1 \mem_reg[20][1]  ( .D(n882), .E(n1008), .CK(clk), .Q(\mem[20][1] ) );
  EDFFX1 \mem_reg[20][0]  ( .D(n876), .E(n1008), .CK(clk), .Q(\mem[20][0] ) );
  EDFFX1 \mem_reg[24][7]  ( .D(n918), .E(n1017), .CK(clk), .Q(\mem[24][7] ) );
  EDFFX1 \mem_reg[24][6]  ( .D(n912), .E(n1017), .CK(clk), .Q(\mem[24][6] ) );
  EDFFX1 \mem_reg[24][5]  ( .D(n906), .E(n1017), .CK(clk), .Q(\mem[24][5] ) );
  EDFFX1 \mem_reg[24][4]  ( .D(n900), .E(n1017), .CK(clk), .Q(\mem[24][4] ) );
  EDFFX1 \mem_reg[24][3]  ( .D(n894), .E(n1017), .CK(clk), .Q(\mem[24][3] ) );
  EDFFX1 \mem_reg[24][2]  ( .D(n888), .E(n1017), .CK(clk), .Q(\mem[24][2] ) );
  EDFFX1 \mem_reg[24][1]  ( .D(n882), .E(n1017), .CK(clk), .Q(\mem[24][1] ) );
  EDFFX1 \mem_reg[24][0]  ( .D(n876), .E(n1017), .CK(clk), .Q(\mem[24][0] ) );
  EDFFX1 \mem_reg[28][7]  ( .D(n918), .E(n1026), .CK(clk), .Q(\mem[28][7] ) );
  EDFFX1 \mem_reg[28][6]  ( .D(n912), .E(n1026), .CK(clk), .Q(\mem[28][6] ) );
  EDFFX1 \mem_reg[28][5]  ( .D(n906), .E(n1026), .CK(clk), .Q(\mem[28][5] ) );
  EDFFX1 \mem_reg[28][4]  ( .D(n900), .E(n1026), .CK(clk), .Q(\mem[28][4] ) );
  EDFFX1 \mem_reg[28][3]  ( .D(n894), .E(n1026), .CK(clk), .Q(\mem[28][3] ) );
  EDFFX1 \mem_reg[28][2]  ( .D(n888), .E(n1026), .CK(clk), .Q(\mem[28][2] ) );
  EDFFX1 \mem_reg[28][1]  ( .D(n882), .E(n1026), .CK(clk), .Q(\mem[28][1] ) );
  EDFFX1 \mem_reg[28][0]  ( .D(n876), .E(n1026), .CK(clk), .Q(\mem[28][0] ) );
  EDFFX1 \mem_reg[32][7]  ( .D(n917), .E(n998), .CK(clk), .Q(\mem[32][7] ) );
  EDFFX1 \mem_reg[32][6]  ( .D(n911), .E(n998), .CK(clk), .Q(\mem[32][6] ) );
  EDFFX1 \mem_reg[32][5]  ( .D(n905), .E(n998), .CK(clk), .Q(\mem[32][5] ) );
  EDFFX1 \mem_reg[32][4]  ( .D(n899), .E(n998), .CK(clk), .Q(\mem[32][4] ) );
  EDFFX1 \mem_reg[32][3]  ( .D(n893), .E(n998), .CK(clk), .Q(\mem[32][3] ) );
  EDFFX1 \mem_reg[32][2]  ( .D(n887), .E(n998), .CK(clk), .Q(\mem[32][2] ) );
  EDFFX1 \mem_reg[32][1]  ( .D(n881), .E(n998), .CK(clk), .Q(\mem[32][1] ) );
  EDFFX1 \mem_reg[32][0]  ( .D(n875), .E(n998), .CK(clk), .Q(\mem[32][0] ) );
  EDFFX1 \mem_reg[36][7]  ( .D(n917), .E(n1007), .CK(clk), .Q(\mem[36][7] ) );
  EDFFX1 \mem_reg[36][6]  ( .D(n911), .E(n1007), .CK(clk), .Q(\mem[36][6] ) );
  EDFFX1 \mem_reg[36][5]  ( .D(n905), .E(n1007), .CK(clk), .Q(\mem[36][5] ) );
  EDFFX1 \mem_reg[36][4]  ( .D(n899), .E(n1007), .CK(clk), .Q(\mem[36][4] ) );
  EDFFX1 \mem_reg[36][3]  ( .D(n893), .E(n1007), .CK(clk), .Q(\mem[36][3] ) );
  EDFFX1 \mem_reg[36][2]  ( .D(n887), .E(n1007), .CK(clk), .Q(\mem[36][2] ) );
  EDFFX1 \mem_reg[36][1]  ( .D(n881), .E(n1007), .CK(clk), .Q(\mem[36][1] ) );
  EDFFX1 \mem_reg[36][0]  ( .D(n875), .E(n1007), .CK(clk), .Q(\mem[36][0] ) );
  EDFFX1 \mem_reg[40][7]  ( .D(n917), .E(n1016), .CK(clk), .Q(\mem[40][7] ) );
  EDFFX1 \mem_reg[40][6]  ( .D(n911), .E(n1016), .CK(clk), .Q(\mem[40][6] ) );
  EDFFX1 \mem_reg[40][5]  ( .D(n905), .E(n1016), .CK(clk), .Q(\mem[40][5] ) );
  EDFFX1 \mem_reg[40][4]  ( .D(n899), .E(n1016), .CK(clk), .Q(\mem[40][4] ) );
  EDFFX1 \mem_reg[40][3]  ( .D(n893), .E(n1016), .CK(clk), .Q(\mem[40][3] ) );
  EDFFX1 \mem_reg[40][2]  ( .D(n887), .E(n1016), .CK(clk), .Q(\mem[40][2] ) );
  EDFFX1 \mem_reg[40][1]  ( .D(n881), .E(n1016), .CK(clk), .Q(\mem[40][1] ) );
  EDFFX1 \mem_reg[40][0]  ( .D(n875), .E(n1016), .CK(clk), .Q(\mem[40][0] ) );
  EDFFX1 \mem_reg[44][7]  ( .D(n916), .E(n1025), .CK(clk), .Q(\mem[44][7] ) );
  EDFFX1 \mem_reg[44][6]  ( .D(n910), .E(n1025), .CK(clk), .Q(\mem[44][6] ) );
  EDFFX1 \mem_reg[44][5]  ( .D(n904), .E(n1025), .CK(clk), .Q(\mem[44][5] ) );
  EDFFX1 \mem_reg[44][4]  ( .D(n898), .E(n1025), .CK(clk), .Q(\mem[44][4] ) );
  EDFFX1 \mem_reg[44][3]  ( .D(n892), .E(n1025), .CK(clk), .Q(\mem[44][3] ) );
  EDFFX1 \mem_reg[44][2]  ( .D(n886), .E(n1025), .CK(clk), .Q(\mem[44][2] ) );
  EDFFX1 \mem_reg[44][1]  ( .D(n880), .E(n1025), .CK(clk), .Q(\mem[44][1] ) );
  EDFFX1 \mem_reg[44][0]  ( .D(n874), .E(n1025), .CK(clk), .Q(\mem[44][0] ) );
  EDFFX1 \mem_reg[48][7]  ( .D(n916), .E(n997), .CK(clk), .Q(\mem[48][7] ) );
  EDFFX1 \mem_reg[48][6]  ( .D(n910), .E(n997), .CK(clk), .Q(\mem[48][6] ) );
  EDFFX1 \mem_reg[48][5]  ( .D(n904), .E(n997), .CK(clk), .Q(\mem[48][5] ) );
  EDFFX1 \mem_reg[48][4]  ( .D(n898), .E(n997), .CK(clk), .Q(\mem[48][4] ) );
  EDFFX1 \mem_reg[48][3]  ( .D(n892), .E(n997), .CK(clk), .Q(\mem[48][3] ) );
  EDFFX1 \mem_reg[48][2]  ( .D(n886), .E(n997), .CK(clk), .Q(\mem[48][2] ) );
  EDFFX1 \mem_reg[48][1]  ( .D(n880), .E(n997), .CK(clk), .Q(\mem[48][1] ) );
  EDFFX1 \mem_reg[48][0]  ( .D(n874), .E(n997), .CK(clk), .Q(\mem[48][0] ) );
  EDFFX1 \mem_reg[52][7]  ( .D(n916), .E(n1006), .CK(clk), .Q(\mem[52][7] ) );
  EDFFX1 \mem_reg[52][6]  ( .D(n910), .E(n1006), .CK(clk), .Q(\mem[52][6] ) );
  EDFFX1 \mem_reg[52][5]  ( .D(n904), .E(n1006), .CK(clk), .Q(\mem[52][5] ) );
  EDFFX1 \mem_reg[52][4]  ( .D(n898), .E(n1006), .CK(clk), .Q(\mem[52][4] ) );
  EDFFX1 \mem_reg[52][3]  ( .D(n892), .E(n1006), .CK(clk), .Q(\mem[52][3] ) );
  EDFFX1 \mem_reg[52][2]  ( .D(n886), .E(n1006), .CK(clk), .Q(\mem[52][2] ) );
  EDFFX1 \mem_reg[52][1]  ( .D(n880), .E(n1006), .CK(clk), .Q(\mem[52][1] ) );
  EDFFX1 \mem_reg[52][0]  ( .D(n874), .E(n1006), .CK(clk), .Q(\mem[52][0] ) );
  EDFFX1 \mem_reg[56][7]  ( .D(n917), .E(n1015), .CK(clk), .Q(\mem[56][7] ) );
  EDFFX1 \mem_reg[56][6]  ( .D(n911), .E(n1015), .CK(clk), .Q(\mem[56][6] ) );
  EDFFX1 \mem_reg[56][5]  ( .D(n905), .E(n1015), .CK(clk), .Q(\mem[56][5] ) );
  EDFFX1 \mem_reg[56][4]  ( .D(n899), .E(n1015), .CK(clk), .Q(\mem[56][4] ) );
  EDFFX1 \mem_reg[56][3]  ( .D(n893), .E(n1015), .CK(clk), .Q(\mem[56][3] ) );
  EDFFX1 \mem_reg[56][2]  ( .D(n887), .E(n1015), .CK(clk), .Q(\mem[56][2] ) );
  EDFFX1 \mem_reg[56][1]  ( .D(n881), .E(n1015), .CK(clk), .Q(\mem[56][1] ) );
  EDFFX1 \mem_reg[56][0]  ( .D(n875), .E(n1015), .CK(clk), .Q(\mem[56][0] ) );
  EDFFX1 \mem_reg[60][7]  ( .D(n914), .E(n1024), .CK(clk), .Q(\mem[60][7] ) );
  EDFFX1 \mem_reg[60][6]  ( .D(n908), .E(n1024), .CK(clk), .Q(\mem[60][6] ) );
  EDFFX1 \mem_reg[60][5]  ( .D(n902), .E(n1024), .CK(clk), .Q(\mem[60][5] ) );
  EDFFX1 \mem_reg[60][4]  ( .D(n896), .E(n1024), .CK(clk), .Q(\mem[60][4] ) );
  EDFFX1 \mem_reg[60][3]  ( .D(n890), .E(n1024), .CK(clk), .Q(\mem[60][3] ) );
  EDFFX1 \mem_reg[60][2]  ( .D(n884), .E(n1024), .CK(clk), .Q(\mem[60][2] ) );
  EDFFX1 \mem_reg[60][1]  ( .D(n878), .E(n1024), .CK(clk), .Q(\mem[60][1] ) );
  EDFFX1 \mem_reg[60][0]  ( .D(n872), .E(n1024), .CK(clk), .Q(\mem[60][0] ) );
  EDFFX1 \mem_reg[64][7]  ( .D(n914), .E(n996), .CK(clk), .Q(\mem[64][7] ) );
  EDFFX1 \mem_reg[64][6]  ( .D(n908), .E(n996), .CK(clk), .Q(\mem[64][6] ) );
  EDFFX1 \mem_reg[64][5]  ( .D(n902), .E(n996), .CK(clk), .Q(\mem[64][5] ) );
  EDFFX1 \mem_reg[64][4]  ( .D(n896), .E(n996), .CK(clk), .Q(\mem[64][4] ) );
  EDFFX1 \mem_reg[64][3]  ( .D(n890), .E(n996), .CK(clk), .Q(\mem[64][3] ) );
  EDFFX1 \mem_reg[64][2]  ( .D(n884), .E(n996), .CK(clk), .Q(\mem[64][2] ) );
  EDFFX1 \mem_reg[64][1]  ( .D(n878), .E(n996), .CK(clk), .Q(\mem[64][1] ) );
  EDFFX1 \mem_reg[64][0]  ( .D(n872), .E(n996), .CK(clk), .Q(\mem[64][0] ) );
  EDFFX1 \mem_reg[68][7]  ( .D(n915), .E(n1005), .CK(clk), .Q(\mem[68][7] ) );
  EDFFX1 \mem_reg[68][6]  ( .D(n909), .E(n1005), .CK(clk), .Q(\mem[68][6] ) );
  EDFFX1 \mem_reg[68][5]  ( .D(n903), .E(n1005), .CK(clk), .Q(\mem[68][5] ) );
  EDFFX1 \mem_reg[68][4]  ( .D(n897), .E(n1005), .CK(clk), .Q(\mem[68][4] ) );
  EDFFX1 \mem_reg[68][3]  ( .D(n891), .E(n1005), .CK(clk), .Q(\mem[68][3] ) );
  EDFFX1 \mem_reg[68][2]  ( .D(n885), .E(n1005), .CK(clk), .Q(\mem[68][2] ) );
  EDFFX1 \mem_reg[68][1]  ( .D(n879), .E(n1005), .CK(clk), .Q(\mem[68][1] ) );
  EDFFX1 \mem_reg[68][0]  ( .D(n873), .E(n1005), .CK(clk), .Q(\mem[68][0] ) );
  EDFFX1 \mem_reg[72][7]  ( .D(n915), .E(n1014), .CK(clk), .Q(\mem[72][7] ) );
  EDFFX1 \mem_reg[72][6]  ( .D(n909), .E(n1014), .CK(clk), .Q(\mem[72][6] ) );
  EDFFX1 \mem_reg[72][5]  ( .D(n903), .E(n1014), .CK(clk), .Q(\mem[72][5] ) );
  EDFFX1 \mem_reg[72][4]  ( .D(n897), .E(n1014), .CK(clk), .Q(\mem[72][4] ) );
  EDFFX1 \mem_reg[72][3]  ( .D(n891), .E(n1014), .CK(clk), .Q(\mem[72][3] ) );
  EDFFX1 \mem_reg[72][2]  ( .D(n885), .E(n1014), .CK(clk), .Q(\mem[72][2] ) );
  EDFFX1 \mem_reg[72][1]  ( .D(n879), .E(n1014), .CK(clk), .Q(\mem[72][1] ) );
  EDFFX1 \mem_reg[72][0]  ( .D(n873), .E(n1014), .CK(clk), .Q(\mem[72][0] ) );
  EDFFX1 \mem_reg[76][7]  ( .D(n915), .E(n1023), .CK(clk), .Q(\mem[76][7] ) );
  EDFFX1 \mem_reg[76][6]  ( .D(n909), .E(n1023), .CK(clk), .Q(\mem[76][6] ) );
  EDFFX1 \mem_reg[76][5]  ( .D(n903), .E(n1023), .CK(clk), .Q(\mem[76][5] ) );
  EDFFX1 \mem_reg[76][4]  ( .D(n897), .E(n1023), .CK(clk), .Q(\mem[76][4] ) );
  EDFFX1 \mem_reg[76][3]  ( .D(n891), .E(n1023), .CK(clk), .Q(\mem[76][3] ) );
  EDFFX1 \mem_reg[76][2]  ( .D(n885), .E(n1023), .CK(clk), .Q(\mem[76][2] ) );
  EDFFX1 \mem_reg[76][1]  ( .D(n879), .E(n1023), .CK(clk), .Q(\mem[76][1] ) );
  EDFFX1 \mem_reg[76][0]  ( .D(n873), .E(n1023), .CK(clk), .Q(\mem[76][0] ) );
  EDFFX1 \mem_reg[80][7]  ( .D(n914), .E(n995), .CK(clk), .Q(\mem[80][7] ) );
  EDFFX1 \mem_reg[80][6]  ( .D(n908), .E(n995), .CK(clk), .Q(\mem[80][6] ) );
  EDFFX1 \mem_reg[80][5]  ( .D(n902), .E(n995), .CK(clk), .Q(\mem[80][5] ) );
  EDFFX1 \mem_reg[80][4]  ( .D(n896), .E(n995), .CK(clk), .Q(\mem[80][4] ) );
  EDFFX1 \mem_reg[80][3]  ( .D(n890), .E(n995), .CK(clk), .Q(\mem[80][3] ) );
  EDFFX1 \mem_reg[80][2]  ( .D(n884), .E(n995), .CK(clk), .Q(\mem[80][2] ) );
  EDFFX1 \mem_reg[80][1]  ( .D(n878), .E(n995), .CK(clk), .Q(\mem[80][1] ) );
  EDFFX1 \mem_reg[80][0]  ( .D(n872), .E(n995), .CK(clk), .Q(\mem[80][0] ) );
  EDFFX1 \mem_reg[84][7]  ( .D(n914), .E(n1004), .CK(clk), .Q(\mem[84][7] ) );
  EDFFX1 \mem_reg[84][6]  ( .D(n908), .E(n1004), .CK(clk), .Q(\mem[84][6] ) );
  EDFFX1 \mem_reg[84][5]  ( .D(n902), .E(n1004), .CK(clk), .Q(\mem[84][5] ) );
  EDFFX1 \mem_reg[84][4]  ( .D(n896), .E(n1004), .CK(clk), .Q(\mem[84][4] ) );
  EDFFX1 \mem_reg[84][3]  ( .D(n890), .E(n1004), .CK(clk), .Q(\mem[84][3] ) );
  EDFFX1 \mem_reg[84][2]  ( .D(n884), .E(n1004), .CK(clk), .Q(\mem[84][2] ) );
  EDFFX1 \mem_reg[84][1]  ( .D(n878), .E(n1004), .CK(clk), .Q(\mem[84][1] ) );
  EDFFX1 \mem_reg[84][0]  ( .D(n872), .E(n1004), .CK(clk), .Q(\mem[84][0] ) );
  EDFFX1 \mem_reg[88][7]  ( .D(n914), .E(n1013), .CK(clk), .Q(\mem[88][7] ) );
  EDFFX1 \mem_reg[88][6]  ( .D(n908), .E(n1013), .CK(clk), .Q(\mem[88][6] ) );
  EDFFX1 \mem_reg[88][5]  ( .D(n902), .E(n1013), .CK(clk), .Q(\mem[88][5] ) );
  EDFFX1 \mem_reg[88][4]  ( .D(n896), .E(n1013), .CK(clk), .Q(\mem[88][4] ) );
  EDFFX1 \mem_reg[88][3]  ( .D(n890), .E(n1013), .CK(clk), .Q(\mem[88][3] ) );
  EDFFX1 \mem_reg[88][2]  ( .D(n884), .E(n1013), .CK(clk), .Q(\mem[88][2] ) );
  EDFFX1 \mem_reg[88][1]  ( .D(n878), .E(n1013), .CK(clk), .Q(\mem[88][1] ) );
  EDFFX1 \mem_reg[88][0]  ( .D(n872), .E(n1013), .CK(clk), .Q(\mem[88][0] ) );
  EDFFX1 \mem_reg[92][7]  ( .D(data_in[7]), .E(n1022), .CK(clk), .Q(
        \mem[92][7] ) );
  EDFFX1 \mem_reg[92][6]  ( .D(data_in[6]), .E(n1022), .CK(clk), .Q(
        \mem[92][6] ) );
  EDFFX1 \mem_reg[92][5]  ( .D(data_in[5]), .E(n1022), .CK(clk), .Q(
        \mem[92][5] ) );
  EDFFX1 \mem_reg[92][4]  ( .D(data_in[4]), .E(n1022), .CK(clk), .Q(
        \mem[92][4] ) );
  EDFFX1 \mem_reg[92][3]  ( .D(data_in[3]), .E(n1022), .CK(clk), .Q(
        \mem[92][3] ) );
  EDFFX1 \mem_reg[92][2]  ( .D(data_in[2]), .E(n1022), .CK(clk), .Q(
        \mem[92][2] ) );
  EDFFX1 \mem_reg[92][1]  ( .D(data_in[1]), .E(n1022), .CK(clk), .Q(
        \mem[92][1] ) );
  EDFFX1 \mem_reg[92][0]  ( .D(data_in[0]), .E(n1022), .CK(clk), .Q(
        \mem[92][0] ) );
  EDFFX1 \mem_reg[96][7]  ( .D(n918), .E(n994), .CK(clk), .Q(\mem[96][7] ) );
  EDFFX1 \mem_reg[96][6]  ( .D(n912), .E(n994), .CK(clk), .Q(\mem[96][6] ) );
  EDFFX1 \mem_reg[96][5]  ( .D(n906), .E(n994), .CK(clk), .Q(\mem[96][5] ) );
  EDFFX1 \mem_reg[96][4]  ( .D(n900), .E(n994), .CK(clk), .Q(\mem[96][4] ) );
  EDFFX1 \mem_reg[96][3]  ( .D(n894), .E(n994), .CK(clk), .Q(\mem[96][3] ) );
  EDFFX1 \mem_reg[96][2]  ( .D(n888), .E(n994), .CK(clk), .Q(\mem[96][2] ) );
  EDFFX1 \mem_reg[96][1]  ( .D(n882), .E(n994), .CK(clk), .Q(\mem[96][1] ) );
  EDFFX1 \mem_reg[96][0]  ( .D(n876), .E(n994), .CK(clk), .Q(\mem[96][0] ) );
  EDFFX1 \mem_reg[100][7]  ( .D(data_in[7]), .E(n1003), .CK(clk), .Q(
        \mem[100][7] ) );
  EDFFX1 \mem_reg[100][6]  ( .D(data_in[6]), .E(n1003), .CK(clk), .Q(
        \mem[100][6] ) );
  EDFFX1 \mem_reg[100][5]  ( .D(data_in[5]), .E(n1003), .CK(clk), .Q(
        \mem[100][5] ) );
  EDFFX1 \mem_reg[100][4]  ( .D(data_in[4]), .E(n1003), .CK(clk), .Q(
        \mem[100][4] ) );
  EDFFX1 \mem_reg[100][3]  ( .D(data_in[3]), .E(n1003), .CK(clk), .Q(
        \mem[100][3] ) );
  EDFFX1 \mem_reg[100][2]  ( .D(data_in[2]), .E(n1003), .CK(clk), .Q(
        \mem[100][2] ) );
  EDFFX1 \mem_reg[100][1]  ( .D(data_in[1]), .E(n1003), .CK(clk), .Q(
        \mem[100][1] ) );
  EDFFX1 \mem_reg[100][0]  ( .D(data_in[0]), .E(n1003), .CK(clk), .Q(
        \mem[100][0] ) );
  EDFFX1 \mem_reg[104][7]  ( .D(n916), .E(n1012), .CK(clk), .Q(\mem[104][7] )
         );
  EDFFX1 \mem_reg[104][6]  ( .D(n910), .E(n1012), .CK(clk), .Q(\mem[104][6] )
         );
  EDFFX1 \mem_reg[104][5]  ( .D(n904), .E(n1012), .CK(clk), .Q(\mem[104][5] )
         );
  EDFFX1 \mem_reg[104][4]  ( .D(n898), .E(n1012), .CK(clk), .Q(\mem[104][4] )
         );
  EDFFX1 \mem_reg[104][3]  ( .D(n892), .E(n1012), .CK(clk), .Q(\mem[104][3] )
         );
  EDFFX1 \mem_reg[104][2]  ( .D(n886), .E(n1012), .CK(clk), .Q(\mem[104][2] )
         );
  EDFFX1 \mem_reg[104][1]  ( .D(n880), .E(n1012), .CK(clk), .Q(\mem[104][1] )
         );
  EDFFX1 \mem_reg[104][0]  ( .D(n874), .E(n1012), .CK(clk), .Q(\mem[104][0] )
         );
  EDFFX1 \mem_reg[108][7]  ( .D(n919), .E(n1021), .CK(clk), .Q(\mem[108][7] )
         );
  EDFFX1 \mem_reg[108][6]  ( .D(n913), .E(n1021), .CK(clk), .Q(\mem[108][6] )
         );
  EDFFX1 \mem_reg[108][5]  ( .D(n907), .E(n1021), .CK(clk), .Q(\mem[108][5] )
         );
  EDFFX1 \mem_reg[108][4]  ( .D(n901), .E(n1021), .CK(clk), .Q(\mem[108][4] )
         );
  EDFFX1 \mem_reg[108][3]  ( .D(n895), .E(n1021), .CK(clk), .Q(\mem[108][3] )
         );
  EDFFX1 \mem_reg[108][2]  ( .D(n889), .E(n1021), .CK(clk), .Q(\mem[108][2] )
         );
  EDFFX1 \mem_reg[108][1]  ( .D(n883), .E(n1021), .CK(clk), .Q(\mem[108][1] )
         );
  EDFFX1 \mem_reg[108][0]  ( .D(n877), .E(n1021), .CK(clk), .Q(\mem[108][0] )
         );
  EDFFX1 \mem_reg[112][7]  ( .D(n917), .E(n993), .CK(clk), .Q(\mem[112][7] )
         );
  EDFFX1 \mem_reg[112][6]  ( .D(n911), .E(n993), .CK(clk), .Q(\mem[112][6] )
         );
  EDFFX1 \mem_reg[112][5]  ( .D(n905), .E(n993), .CK(clk), .Q(\mem[112][5] )
         );
  EDFFX1 \mem_reg[112][4]  ( .D(n899), .E(n993), .CK(clk), .Q(\mem[112][4] )
         );
  EDFFX1 \mem_reg[112][3]  ( .D(n893), .E(n993), .CK(clk), .Q(\mem[112][3] )
         );
  EDFFX1 \mem_reg[112][2]  ( .D(n887), .E(n993), .CK(clk), .Q(\mem[112][2] )
         );
  EDFFX1 \mem_reg[112][1]  ( .D(n881), .E(n993), .CK(clk), .Q(\mem[112][1] )
         );
  EDFFX1 \mem_reg[112][0]  ( .D(n875), .E(n993), .CK(clk), .Q(\mem[112][0] )
         );
  EDFFX1 \mem_reg[116][7]  ( .D(n918), .E(n1002), .CK(clk), .Q(\mem[116][7] )
         );
  EDFFX1 \mem_reg[116][6]  ( .D(n912), .E(n1002), .CK(clk), .Q(\mem[116][6] )
         );
  EDFFX1 \mem_reg[116][5]  ( .D(n906), .E(n1002), .CK(clk), .Q(\mem[116][5] )
         );
  EDFFX1 \mem_reg[116][4]  ( .D(n900), .E(n1002), .CK(clk), .Q(\mem[116][4] )
         );
  EDFFX1 \mem_reg[116][3]  ( .D(n894), .E(n1002), .CK(clk), .Q(\mem[116][3] )
         );
  EDFFX1 \mem_reg[116][2]  ( .D(n888), .E(n1002), .CK(clk), .Q(\mem[116][2] )
         );
  EDFFX1 \mem_reg[116][1]  ( .D(n882), .E(n1002), .CK(clk), .Q(\mem[116][1] )
         );
  EDFFX1 \mem_reg[116][0]  ( .D(n876), .E(n1002), .CK(clk), .Q(\mem[116][0] )
         );
  EDFFX1 \mem_reg[120][7]  ( .D(n916), .E(n1011), .CK(clk), .Q(\mem[120][7] )
         );
  EDFFX1 \mem_reg[120][6]  ( .D(n910), .E(n1011), .CK(clk), .Q(\mem[120][6] )
         );
  EDFFX1 \mem_reg[120][5]  ( .D(n904), .E(n1011), .CK(clk), .Q(\mem[120][5] )
         );
  EDFFX1 \mem_reg[120][4]  ( .D(n898), .E(n1011), .CK(clk), .Q(\mem[120][4] )
         );
  EDFFX1 \mem_reg[120][3]  ( .D(n892), .E(n1011), .CK(clk), .Q(\mem[120][3] )
         );
  EDFFX1 \mem_reg[120][2]  ( .D(n886), .E(n1011), .CK(clk), .Q(\mem[120][2] )
         );
  EDFFX1 \mem_reg[120][1]  ( .D(n880), .E(n1011), .CK(clk), .Q(\mem[120][1] )
         );
  EDFFX1 \mem_reg[120][0]  ( .D(n874), .E(n1011), .CK(clk), .Q(\mem[120][0] )
         );
  EDFFX1 \mem_reg[124][7]  ( .D(n919), .E(n1020), .CK(clk), .Q(\mem[124][7] )
         );
  EDFFX1 \mem_reg[124][6]  ( .D(n913), .E(n1020), .CK(clk), .Q(\mem[124][6] )
         );
  EDFFX1 \mem_reg[124][5]  ( .D(n907), .E(n1020), .CK(clk), .Q(\mem[124][5] )
         );
  EDFFX1 \mem_reg[124][4]  ( .D(n901), .E(n1020), .CK(clk), .Q(\mem[124][4] )
         );
  EDFFX1 \mem_reg[124][3]  ( .D(n895), .E(n1020), .CK(clk), .Q(\mem[124][3] )
         );
  EDFFX1 \mem_reg[124][2]  ( .D(n889), .E(n1020), .CK(clk), .Q(\mem[124][2] )
         );
  EDFFX1 \mem_reg[124][1]  ( .D(n883), .E(n1020), .CK(clk), .Q(\mem[124][1] )
         );
  EDFFX1 \mem_reg[124][0]  ( .D(n877), .E(n1020), .CK(clk), .Q(\mem[124][0] )
         );
  EDFFX1 \mem_reg[2][7]  ( .D(n915), .E(n1036), .CK(clk), .Q(\mem[2][7] ) );
  EDFFX1 \mem_reg[2][6]  ( .D(n909), .E(n1036), .CK(clk), .Q(\mem[2][6] ) );
  EDFFX1 \mem_reg[2][5]  ( .D(n903), .E(n1036), .CK(clk), .Q(\mem[2][5] ) );
  EDFFX1 \mem_reg[2][4]  ( .D(n897), .E(n1036), .CK(clk), .Q(\mem[2][4] ) );
  EDFFX1 \mem_reg[2][3]  ( .D(n891), .E(n1036), .CK(clk), .Q(\mem[2][3] ) );
  EDFFX1 \mem_reg[2][2]  ( .D(n885), .E(n1036), .CK(clk), .Q(\mem[2][2] ) );
  EDFFX1 \mem_reg[2][1]  ( .D(n879), .E(n1036), .CK(clk), .Q(\mem[2][1] ) );
  EDFFX1 \mem_reg[2][0]  ( .D(n873), .E(n1036), .CK(clk), .Q(\mem[2][0] ) );
  EDFFX1 \mem_reg[6][7]  ( .D(n914), .E(n1045), .CK(clk), .Q(\mem[6][7] ) );
  EDFFX1 \mem_reg[6][6]  ( .D(n908), .E(n1045), .CK(clk), .Q(\mem[6][6] ) );
  EDFFX1 \mem_reg[6][5]  ( .D(n902), .E(n1045), .CK(clk), .Q(\mem[6][5] ) );
  EDFFX1 \mem_reg[6][4]  ( .D(n896), .E(n1045), .CK(clk), .Q(\mem[6][4] ) );
  EDFFX1 \mem_reg[6][3]  ( .D(n890), .E(n1045), .CK(clk), .Q(\mem[6][3] ) );
  EDFFX1 \mem_reg[6][2]  ( .D(n884), .E(n1045), .CK(clk), .Q(\mem[6][2] ) );
  EDFFX1 \mem_reg[6][1]  ( .D(n878), .E(n1045), .CK(clk), .Q(\mem[6][1] ) );
  EDFFX1 \mem_reg[6][0]  ( .D(n872), .E(n1045), .CK(clk), .Q(\mem[6][0] ) );
  EDFFX1 \mem_reg[10][7]  ( .D(n919), .E(n1054), .CK(clk), .Q(\mem[10][7] ) );
  EDFFX1 \mem_reg[10][6]  ( .D(n913), .E(n1054), .CK(clk), .Q(\mem[10][6] ) );
  EDFFX1 \mem_reg[10][5]  ( .D(n907), .E(n1054), .CK(clk), .Q(\mem[10][5] ) );
  EDFFX1 \mem_reg[10][4]  ( .D(n901), .E(n1054), .CK(clk), .Q(\mem[10][4] ) );
  EDFFX1 \mem_reg[10][3]  ( .D(n895), .E(n1054), .CK(clk), .Q(\mem[10][3] ) );
  EDFFX1 \mem_reg[10][2]  ( .D(n889), .E(n1054), .CK(clk), .Q(\mem[10][2] ) );
  EDFFX1 \mem_reg[10][1]  ( .D(n883), .E(n1054), .CK(clk), .Q(\mem[10][1] ) );
  EDFFX1 \mem_reg[10][0]  ( .D(n877), .E(n1054), .CK(clk), .Q(\mem[10][0] ) );
  EDFFX1 \mem_reg[14][7]  ( .D(n919), .E(n1063), .CK(clk), .Q(\mem[14][7] ) );
  EDFFX1 \mem_reg[14][6]  ( .D(n913), .E(n1063), .CK(clk), .Q(\mem[14][6] ) );
  EDFFX1 \mem_reg[14][5]  ( .D(n907), .E(n1063), .CK(clk), .Q(\mem[14][5] ) );
  EDFFX1 \mem_reg[14][4]  ( .D(n901), .E(n1063), .CK(clk), .Q(\mem[14][4] ) );
  EDFFX1 \mem_reg[14][3]  ( .D(n895), .E(n1063), .CK(clk), .Q(\mem[14][3] ) );
  EDFFX1 \mem_reg[14][2]  ( .D(n889), .E(n1063), .CK(clk), .Q(\mem[14][2] ) );
  EDFFX1 \mem_reg[14][1]  ( .D(n883), .E(n1063), .CK(clk), .Q(\mem[14][1] ) );
  EDFFX1 \mem_reg[14][0]  ( .D(n877), .E(n1063), .CK(clk), .Q(\mem[14][0] ) );
  EDFFX1 \mem_reg[18][7]  ( .D(n919), .E(n1035), .CK(clk), .Q(\mem[18][7] ) );
  EDFFX1 \mem_reg[18][6]  ( .D(n913), .E(n1035), .CK(clk), .Q(\mem[18][6] ) );
  EDFFX1 \mem_reg[18][5]  ( .D(n907), .E(n1035), .CK(clk), .Q(\mem[18][5] ) );
  EDFFX1 \mem_reg[18][4]  ( .D(n901), .E(n1035), .CK(clk), .Q(\mem[18][4] ) );
  EDFFX1 \mem_reg[18][3]  ( .D(n895), .E(n1035), .CK(clk), .Q(\mem[18][3] ) );
  EDFFX1 \mem_reg[18][2]  ( .D(n889), .E(n1035), .CK(clk), .Q(\mem[18][2] ) );
  EDFFX1 \mem_reg[18][1]  ( .D(n883), .E(n1035), .CK(clk), .Q(\mem[18][1] ) );
  EDFFX1 \mem_reg[18][0]  ( .D(n877), .E(n1035), .CK(clk), .Q(\mem[18][0] ) );
  EDFFX1 \mem_reg[22][7]  ( .D(n918), .E(n1044), .CK(clk), .Q(\mem[22][7] ) );
  EDFFX1 \mem_reg[22][6]  ( .D(n912), .E(n1044), .CK(clk), .Q(\mem[22][6] ) );
  EDFFX1 \mem_reg[22][5]  ( .D(n906), .E(n1044), .CK(clk), .Q(\mem[22][5] ) );
  EDFFX1 \mem_reg[22][4]  ( .D(n900), .E(n1044), .CK(clk), .Q(\mem[22][4] ) );
  EDFFX1 \mem_reg[22][3]  ( .D(n894), .E(n1044), .CK(clk), .Q(\mem[22][3] ) );
  EDFFX1 \mem_reg[22][2]  ( .D(n888), .E(n1044), .CK(clk), .Q(\mem[22][2] ) );
  EDFFX1 \mem_reg[22][1]  ( .D(n882), .E(n1044), .CK(clk), .Q(\mem[22][1] ) );
  EDFFX1 \mem_reg[22][0]  ( .D(n876), .E(n1044), .CK(clk), .Q(\mem[22][0] ) );
  EDFFX1 \mem_reg[26][7]  ( .D(n918), .E(n1053), .CK(clk), .Q(\mem[26][7] ) );
  EDFFX1 \mem_reg[26][6]  ( .D(n912), .E(n1053), .CK(clk), .Q(\mem[26][6] ) );
  EDFFX1 \mem_reg[26][5]  ( .D(n906), .E(n1053), .CK(clk), .Q(\mem[26][5] ) );
  EDFFX1 \mem_reg[26][4]  ( .D(n900), .E(n1053), .CK(clk), .Q(\mem[26][4] ) );
  EDFFX1 \mem_reg[26][3]  ( .D(n894), .E(n1053), .CK(clk), .Q(\mem[26][3] ) );
  EDFFX1 \mem_reg[26][2]  ( .D(n888), .E(n1053), .CK(clk), .Q(\mem[26][2] ) );
  EDFFX1 \mem_reg[26][1]  ( .D(n882), .E(n1053), .CK(clk), .Q(\mem[26][1] ) );
  EDFFX1 \mem_reg[26][0]  ( .D(n876), .E(n1053), .CK(clk), .Q(\mem[26][0] ) );
  EDFFX1 \mem_reg[30][7]  ( .D(n918), .E(n1062), .CK(clk), .Q(\mem[30][7] ) );
  EDFFX1 \mem_reg[30][6]  ( .D(n912), .E(n1062), .CK(clk), .Q(\mem[30][6] ) );
  EDFFX1 \mem_reg[30][5]  ( .D(n906), .E(n1062), .CK(clk), .Q(\mem[30][5] ) );
  EDFFX1 \mem_reg[30][4]  ( .D(n900), .E(n1062), .CK(clk), .Q(\mem[30][4] ) );
  EDFFX1 \mem_reg[30][3]  ( .D(n894), .E(n1062), .CK(clk), .Q(\mem[30][3] ) );
  EDFFX1 \mem_reg[30][2]  ( .D(n888), .E(n1062), .CK(clk), .Q(\mem[30][2] ) );
  EDFFX1 \mem_reg[30][1]  ( .D(n882), .E(n1062), .CK(clk), .Q(\mem[30][1] ) );
  EDFFX1 \mem_reg[30][0]  ( .D(n876), .E(n1062), .CK(clk), .Q(\mem[30][0] ) );
  EDFFX1 \mem_reg[34][7]  ( .D(n917), .E(n1034), .CK(clk), .Q(\mem[34][7] ) );
  EDFFX1 \mem_reg[34][6]  ( .D(n911), .E(n1034), .CK(clk), .Q(\mem[34][6] ) );
  EDFFX1 \mem_reg[34][5]  ( .D(n905), .E(n1034), .CK(clk), .Q(\mem[34][5] ) );
  EDFFX1 \mem_reg[34][4]  ( .D(n899), .E(n1034), .CK(clk), .Q(\mem[34][4] ) );
  EDFFX1 \mem_reg[34][3]  ( .D(n893), .E(n1034), .CK(clk), .Q(\mem[34][3] ) );
  EDFFX1 \mem_reg[34][2]  ( .D(n887), .E(n1034), .CK(clk), .Q(\mem[34][2] ) );
  EDFFX1 \mem_reg[34][1]  ( .D(n881), .E(n1034), .CK(clk), .Q(\mem[34][1] ) );
  EDFFX1 \mem_reg[34][0]  ( .D(n875), .E(n1034), .CK(clk), .Q(\mem[34][0] ) );
  EDFFX1 \mem_reg[38][7]  ( .D(n917), .E(n1043), .CK(clk), .Q(\mem[38][7] ) );
  EDFFX1 \mem_reg[38][6]  ( .D(n911), .E(n1043), .CK(clk), .Q(\mem[38][6] ) );
  EDFFX1 \mem_reg[38][5]  ( .D(n905), .E(n1043), .CK(clk), .Q(\mem[38][5] ) );
  EDFFX1 \mem_reg[38][4]  ( .D(n899), .E(n1043), .CK(clk), .Q(\mem[38][4] ) );
  EDFFX1 \mem_reg[38][3]  ( .D(n893), .E(n1043), .CK(clk), .Q(\mem[38][3] ) );
  EDFFX1 \mem_reg[38][2]  ( .D(n887), .E(n1043), .CK(clk), .Q(\mem[38][2] ) );
  EDFFX1 \mem_reg[38][1]  ( .D(n881), .E(n1043), .CK(clk), .Q(\mem[38][1] ) );
  EDFFX1 \mem_reg[38][0]  ( .D(n875), .E(n1043), .CK(clk), .Q(\mem[38][0] ) );
  EDFFX1 \mem_reg[42][7]  ( .D(n917), .E(n1052), .CK(clk), .Q(\mem[42][7] ) );
  EDFFX1 \mem_reg[42][6]  ( .D(n911), .E(n1052), .CK(clk), .Q(\mem[42][6] ) );
  EDFFX1 \mem_reg[42][5]  ( .D(n905), .E(n1052), .CK(clk), .Q(\mem[42][5] ) );
  EDFFX1 \mem_reg[42][4]  ( .D(n899), .E(n1052), .CK(clk), .Q(\mem[42][4] ) );
  EDFFX1 \mem_reg[42][3]  ( .D(n893), .E(n1052), .CK(clk), .Q(\mem[42][3] ) );
  EDFFX1 \mem_reg[42][2]  ( .D(n887), .E(n1052), .CK(clk), .Q(\mem[42][2] ) );
  EDFFX1 \mem_reg[42][1]  ( .D(n881), .E(n1052), .CK(clk), .Q(\mem[42][1] ) );
  EDFFX1 \mem_reg[42][0]  ( .D(n875), .E(n1052), .CK(clk), .Q(\mem[42][0] ) );
  EDFFX1 \mem_reg[46][7]  ( .D(n916), .E(n1061), .CK(clk), .Q(\mem[46][7] ) );
  EDFFX1 \mem_reg[46][6]  ( .D(n910), .E(n1061), .CK(clk), .Q(\mem[46][6] ) );
  EDFFX1 \mem_reg[46][5]  ( .D(n904), .E(n1061), .CK(clk), .Q(\mem[46][5] ) );
  EDFFX1 \mem_reg[46][4]  ( .D(n898), .E(n1061), .CK(clk), .Q(\mem[46][4] ) );
  EDFFX1 \mem_reg[46][3]  ( .D(n892), .E(n1061), .CK(clk), .Q(\mem[46][3] ) );
  EDFFX1 \mem_reg[46][2]  ( .D(n886), .E(n1061), .CK(clk), .Q(\mem[46][2] ) );
  EDFFX1 \mem_reg[46][1]  ( .D(n880), .E(n1061), .CK(clk), .Q(\mem[46][1] ) );
  EDFFX1 \mem_reg[46][0]  ( .D(n874), .E(n1061), .CK(clk), .Q(\mem[46][0] ) );
  EDFFX1 \mem_reg[50][7]  ( .D(n916), .E(n1033), .CK(clk), .Q(\mem[50][7] ) );
  EDFFX1 \mem_reg[50][6]  ( .D(n910), .E(n1033), .CK(clk), .Q(\mem[50][6] ) );
  EDFFX1 \mem_reg[50][5]  ( .D(n904), .E(n1033), .CK(clk), .Q(\mem[50][5] ) );
  EDFFX1 \mem_reg[50][4]  ( .D(n898), .E(n1033), .CK(clk), .Q(\mem[50][4] ) );
  EDFFX1 \mem_reg[50][3]  ( .D(n892), .E(n1033), .CK(clk), .Q(\mem[50][3] ) );
  EDFFX1 \mem_reg[50][2]  ( .D(n886), .E(n1033), .CK(clk), .Q(\mem[50][2] ) );
  EDFFX1 \mem_reg[50][1]  ( .D(n880), .E(n1033), .CK(clk), .Q(\mem[50][1] ) );
  EDFFX1 \mem_reg[50][0]  ( .D(n874), .E(n1033), .CK(clk), .Q(\mem[50][0] ) );
  EDFFX1 \mem_reg[54][7]  ( .D(n916), .E(n1042), .CK(clk), .Q(\mem[54][7] ) );
  EDFFX1 \mem_reg[54][6]  ( .D(n910), .E(n1042), .CK(clk), .Q(\mem[54][6] ) );
  EDFFX1 \mem_reg[54][5]  ( .D(n904), .E(n1042), .CK(clk), .Q(\mem[54][5] ) );
  EDFFX1 \mem_reg[54][4]  ( .D(n898), .E(n1042), .CK(clk), .Q(\mem[54][4] ) );
  EDFFX1 \mem_reg[54][3]  ( .D(n892), .E(n1042), .CK(clk), .Q(\mem[54][3] ) );
  EDFFX1 \mem_reg[54][2]  ( .D(n886), .E(n1042), .CK(clk), .Q(\mem[54][2] ) );
  EDFFX1 \mem_reg[54][1]  ( .D(n880), .E(n1042), .CK(clk), .Q(\mem[54][1] ) );
  EDFFX1 \mem_reg[54][0]  ( .D(n874), .E(n1042), .CK(clk), .Q(\mem[54][0] ) );
  EDFFX1 \mem_reg[58][7]  ( .D(n915), .E(n1051), .CK(clk), .Q(\mem[58][7] ) );
  EDFFX1 \mem_reg[58][6]  ( .D(n909), .E(n1051), .CK(clk), .Q(\mem[58][6] ) );
  EDFFX1 \mem_reg[58][5]  ( .D(n903), .E(n1051), .CK(clk), .Q(\mem[58][5] ) );
  EDFFX1 \mem_reg[58][4]  ( .D(n897), .E(n1051), .CK(clk), .Q(\mem[58][4] ) );
  EDFFX1 \mem_reg[58][3]  ( .D(n891), .E(n1051), .CK(clk), .Q(\mem[58][3] ) );
  EDFFX1 \mem_reg[58][2]  ( .D(n885), .E(n1051), .CK(clk), .Q(\mem[58][2] ) );
  EDFFX1 \mem_reg[58][1]  ( .D(n879), .E(n1051), .CK(clk), .Q(\mem[58][1] ) );
  EDFFX1 \mem_reg[58][0]  ( .D(n873), .E(n1051), .CK(clk), .Q(\mem[58][0] ) );
  EDFFX1 \mem_reg[62][7]  ( .D(n918), .E(n1060), .CK(clk), .Q(\mem[62][7] ) );
  EDFFX1 \mem_reg[62][6]  ( .D(n912), .E(n1060), .CK(clk), .Q(\mem[62][6] ) );
  EDFFX1 \mem_reg[62][5]  ( .D(n906), .E(n1060), .CK(clk), .Q(\mem[62][5] ) );
  EDFFX1 \mem_reg[62][4]  ( .D(n900), .E(n1060), .CK(clk), .Q(\mem[62][4] ) );
  EDFFX1 \mem_reg[62][3]  ( .D(n894), .E(n1060), .CK(clk), .Q(\mem[62][3] ) );
  EDFFX1 \mem_reg[62][2]  ( .D(n888), .E(n1060), .CK(clk), .Q(\mem[62][2] ) );
  EDFFX1 \mem_reg[62][1]  ( .D(n882), .E(n1060), .CK(clk), .Q(\mem[62][1] ) );
  EDFFX1 \mem_reg[62][0]  ( .D(n876), .E(n1060), .CK(clk), .Q(\mem[62][0] ) );
  EDFFX1 \mem_reg[66][7]  ( .D(data_in[7]), .E(n1032), .CK(clk), .Q(
        \mem[66][7] ) );
  EDFFX1 \mem_reg[66][6]  ( .D(data_in[6]), .E(n1032), .CK(clk), .Q(
        \mem[66][6] ) );
  EDFFX1 \mem_reg[66][5]  ( .D(data_in[5]), .E(n1032), .CK(clk), .Q(
        \mem[66][5] ) );
  EDFFX1 \mem_reg[66][4]  ( .D(data_in[4]), .E(n1032), .CK(clk), .Q(
        \mem[66][4] ) );
  EDFFX1 \mem_reg[66][3]  ( .D(data_in[3]), .E(n1032), .CK(clk), .Q(
        \mem[66][3] ) );
  EDFFX1 \mem_reg[66][2]  ( .D(data_in[2]), .E(n1032), .CK(clk), .Q(
        \mem[66][2] ) );
  EDFFX1 \mem_reg[66][1]  ( .D(data_in[1]), .E(n1032), .CK(clk), .Q(
        \mem[66][1] ) );
  EDFFX1 \mem_reg[66][0]  ( .D(data_in[0]), .E(n1032), .CK(clk), .Q(
        \mem[66][0] ) );
  EDFFX1 \mem_reg[70][7]  ( .D(n915), .E(n1041), .CK(clk), .Q(\mem[70][7] ) );
  EDFFX1 \mem_reg[70][6]  ( .D(n909), .E(n1041), .CK(clk), .Q(\mem[70][6] ) );
  EDFFX1 \mem_reg[70][5]  ( .D(n903), .E(n1041), .CK(clk), .Q(\mem[70][5] ) );
  EDFFX1 \mem_reg[70][4]  ( .D(n897), .E(n1041), .CK(clk), .Q(\mem[70][4] ) );
  EDFFX1 \mem_reg[70][3]  ( .D(n891), .E(n1041), .CK(clk), .Q(\mem[70][3] ) );
  EDFFX1 \mem_reg[70][2]  ( .D(n885), .E(n1041), .CK(clk), .Q(\mem[70][2] ) );
  EDFFX1 \mem_reg[70][1]  ( .D(n879), .E(n1041), .CK(clk), .Q(\mem[70][1] ) );
  EDFFX1 \mem_reg[70][0]  ( .D(n873), .E(n1041), .CK(clk), .Q(\mem[70][0] ) );
  EDFFX1 \mem_reg[74][7]  ( .D(n915), .E(n1050), .CK(clk), .Q(\mem[74][7] ) );
  EDFFX1 \mem_reg[74][6]  ( .D(n909), .E(n1050), .CK(clk), .Q(\mem[74][6] ) );
  EDFFX1 \mem_reg[74][5]  ( .D(n903), .E(n1050), .CK(clk), .Q(\mem[74][5] ) );
  EDFFX1 \mem_reg[74][4]  ( .D(n897), .E(n1050), .CK(clk), .Q(\mem[74][4] ) );
  EDFFX1 \mem_reg[74][3]  ( .D(n891), .E(n1050), .CK(clk), .Q(\mem[74][3] ) );
  EDFFX1 \mem_reg[74][2]  ( .D(n885), .E(n1050), .CK(clk), .Q(\mem[74][2] ) );
  EDFFX1 \mem_reg[74][1]  ( .D(n879), .E(n1050), .CK(clk), .Q(\mem[74][1] ) );
  EDFFX1 \mem_reg[74][0]  ( .D(n873), .E(n1050), .CK(clk), .Q(\mem[74][0] ) );
  EDFFX1 \mem_reg[78][7]  ( .D(n915), .E(n1059), .CK(clk), .Q(\mem[78][7] ) );
  EDFFX1 \mem_reg[78][6]  ( .D(n909), .E(n1059), .CK(clk), .Q(\mem[78][6] ) );
  EDFFX1 \mem_reg[78][5]  ( .D(n903), .E(n1059), .CK(clk), .Q(\mem[78][5] ) );
  EDFFX1 \mem_reg[78][4]  ( .D(n897), .E(n1059), .CK(clk), .Q(\mem[78][4] ) );
  EDFFX1 \mem_reg[78][3]  ( .D(n891), .E(n1059), .CK(clk), .Q(\mem[78][3] ) );
  EDFFX1 \mem_reg[78][2]  ( .D(n885), .E(n1059), .CK(clk), .Q(\mem[78][2] ) );
  EDFFX1 \mem_reg[78][1]  ( .D(n879), .E(n1059), .CK(clk), .Q(\mem[78][1] ) );
  EDFFX1 \mem_reg[78][0]  ( .D(n873), .E(n1059), .CK(clk), .Q(\mem[78][0] ) );
  EDFFX1 \mem_reg[82][7]  ( .D(n914), .E(n1031), .CK(clk), .Q(\mem[82][7] ) );
  EDFFX1 \mem_reg[82][6]  ( .D(n908), .E(n1031), .CK(clk), .Q(\mem[82][6] ) );
  EDFFX1 \mem_reg[82][5]  ( .D(n902), .E(n1031), .CK(clk), .Q(\mem[82][5] ) );
  EDFFX1 \mem_reg[82][4]  ( .D(n896), .E(n1031), .CK(clk), .Q(\mem[82][4] ) );
  EDFFX1 \mem_reg[82][3]  ( .D(n890), .E(n1031), .CK(clk), .Q(\mem[82][3] ) );
  EDFFX1 \mem_reg[82][2]  ( .D(n884), .E(n1031), .CK(clk), .Q(\mem[82][2] ) );
  EDFFX1 \mem_reg[82][1]  ( .D(n878), .E(n1031), .CK(clk), .Q(\mem[82][1] ) );
  EDFFX1 \mem_reg[82][0]  ( .D(n872), .E(n1031), .CK(clk), .Q(\mem[82][0] ) );
  EDFFX1 \mem_reg[86][7]  ( .D(n914), .E(n1040), .CK(clk), .Q(\mem[86][7] ) );
  EDFFX1 \mem_reg[86][6]  ( .D(n908), .E(n1040), .CK(clk), .Q(\mem[86][6] ) );
  EDFFX1 \mem_reg[86][5]  ( .D(n902), .E(n1040), .CK(clk), .Q(\mem[86][5] ) );
  EDFFX1 \mem_reg[86][4]  ( .D(n896), .E(n1040), .CK(clk), .Q(\mem[86][4] ) );
  EDFFX1 \mem_reg[86][3]  ( .D(n890), .E(n1040), .CK(clk), .Q(\mem[86][3] ) );
  EDFFX1 \mem_reg[86][2]  ( .D(n884), .E(n1040), .CK(clk), .Q(\mem[86][2] ) );
  EDFFX1 \mem_reg[86][1]  ( .D(n878), .E(n1040), .CK(clk), .Q(\mem[86][1] ) );
  EDFFX1 \mem_reg[86][0]  ( .D(n872), .E(n1040), .CK(clk), .Q(\mem[86][0] ) );
  EDFFX1 \mem_reg[90][7]  ( .D(n914), .E(n1049), .CK(clk), .Q(\mem[90][7] ) );
  EDFFX1 \mem_reg[90][6]  ( .D(n908), .E(n1049), .CK(clk), .Q(\mem[90][6] ) );
  EDFFX1 \mem_reg[90][5]  ( .D(n902), .E(n1049), .CK(clk), .Q(\mem[90][5] ) );
  EDFFX1 \mem_reg[90][4]  ( .D(n896), .E(n1049), .CK(clk), .Q(\mem[90][4] ) );
  EDFFX1 \mem_reg[90][3]  ( .D(n890), .E(n1049), .CK(clk), .Q(\mem[90][3] ) );
  EDFFX1 \mem_reg[90][2]  ( .D(n884), .E(n1049), .CK(clk), .Q(\mem[90][2] ) );
  EDFFX1 \mem_reg[90][1]  ( .D(n878), .E(n1049), .CK(clk), .Q(\mem[90][1] ) );
  EDFFX1 \mem_reg[90][0]  ( .D(n872), .E(n1049), .CK(clk), .Q(\mem[90][0] ) );
  EDFFX1 \mem_reg[94][7]  ( .D(n916), .E(n1058), .CK(clk), .Q(\mem[94][7] ) );
  EDFFX1 \mem_reg[94][6]  ( .D(n910), .E(n1058), .CK(clk), .Q(\mem[94][6] ) );
  EDFFX1 \mem_reg[94][5]  ( .D(n904), .E(n1058), .CK(clk), .Q(\mem[94][5] ) );
  EDFFX1 \mem_reg[94][4]  ( .D(n898), .E(n1058), .CK(clk), .Q(\mem[94][4] ) );
  EDFFX1 \mem_reg[94][3]  ( .D(n892), .E(n1058), .CK(clk), .Q(\mem[94][3] ) );
  EDFFX1 \mem_reg[94][2]  ( .D(n886), .E(n1058), .CK(clk), .Q(\mem[94][2] ) );
  EDFFX1 \mem_reg[94][1]  ( .D(n880), .E(n1058), .CK(clk), .Q(\mem[94][1] ) );
  EDFFX1 \mem_reg[94][0]  ( .D(n874), .E(n1058), .CK(clk), .Q(\mem[94][0] ) );
  EDFFX1 \mem_reg[98][7]  ( .D(data_in[7]), .E(n1030), .CK(clk), .Q(
        \mem[98][7] ) );
  EDFFX1 \mem_reg[98][6]  ( .D(data_in[6]), .E(n1030), .CK(clk), .Q(
        \mem[98][6] ) );
  EDFFX1 \mem_reg[98][5]  ( .D(data_in[5]), .E(n1030), .CK(clk), .Q(
        \mem[98][5] ) );
  EDFFX1 \mem_reg[98][4]  ( .D(data_in[4]), .E(n1030), .CK(clk), .Q(
        \mem[98][4] ) );
  EDFFX1 \mem_reg[98][3]  ( .D(data_in[3]), .E(n1030), .CK(clk), .Q(
        \mem[98][3] ) );
  EDFFX1 \mem_reg[98][2]  ( .D(data_in[2]), .E(n1030), .CK(clk), .Q(
        \mem[98][2] ) );
  EDFFX1 \mem_reg[98][1]  ( .D(data_in[1]), .E(n1030), .CK(clk), .Q(
        \mem[98][1] ) );
  EDFFX1 \mem_reg[98][0]  ( .D(data_in[0]), .E(n1030), .CK(clk), .Q(
        \mem[98][0] ) );
  EDFFX1 \mem_reg[102][7]  ( .D(n919), .E(n1039), .CK(clk), .Q(\mem[102][7] )
         );
  EDFFX1 \mem_reg[102][6]  ( .D(n913), .E(n1039), .CK(clk), .Q(\mem[102][6] )
         );
  EDFFX1 \mem_reg[102][5]  ( .D(n907), .E(n1039), .CK(clk), .Q(\mem[102][5] )
         );
  EDFFX1 \mem_reg[102][4]  ( .D(n901), .E(n1039), .CK(clk), .Q(\mem[102][4] )
         );
  EDFFX1 \mem_reg[102][3]  ( .D(n895), .E(n1039), .CK(clk), .Q(\mem[102][3] )
         );
  EDFFX1 \mem_reg[102][2]  ( .D(n889), .E(n1039), .CK(clk), .Q(\mem[102][2] )
         );
  EDFFX1 \mem_reg[102][1]  ( .D(n883), .E(n1039), .CK(clk), .Q(\mem[102][1] )
         );
  EDFFX1 \mem_reg[102][0]  ( .D(n877), .E(n1039), .CK(clk), .Q(\mem[102][0] )
         );
  EDFFX1 \mem_reg[106][7]  ( .D(n917), .E(n1048), .CK(clk), .Q(\mem[106][7] )
         );
  EDFFX1 \mem_reg[106][6]  ( .D(n911), .E(n1048), .CK(clk), .Q(\mem[106][6] )
         );
  EDFFX1 \mem_reg[106][5]  ( .D(n905), .E(n1048), .CK(clk), .Q(\mem[106][5] )
         );
  EDFFX1 \mem_reg[106][4]  ( .D(n899), .E(n1048), .CK(clk), .Q(\mem[106][4] )
         );
  EDFFX1 \mem_reg[106][3]  ( .D(n893), .E(n1048), .CK(clk), .Q(\mem[106][3] )
         );
  EDFFX1 \mem_reg[106][2]  ( .D(n887), .E(n1048), .CK(clk), .Q(\mem[106][2] )
         );
  EDFFX1 \mem_reg[106][1]  ( .D(n881), .E(n1048), .CK(clk), .Q(\mem[106][1] )
         );
  EDFFX1 \mem_reg[106][0]  ( .D(n875), .E(n1048), .CK(clk), .Q(\mem[106][0] )
         );
  EDFFX1 \mem_reg[110][7]  ( .D(n918), .E(n1057), .CK(clk), .Q(\mem[110][7] )
         );
  EDFFX1 \mem_reg[110][6]  ( .D(n912), .E(n1057), .CK(clk), .Q(\mem[110][6] )
         );
  EDFFX1 \mem_reg[110][5]  ( .D(n906), .E(n1057), .CK(clk), .Q(\mem[110][5] )
         );
  EDFFX1 \mem_reg[110][4]  ( .D(n900), .E(n1057), .CK(clk), .Q(\mem[110][4] )
         );
  EDFFX1 \mem_reg[110][3]  ( .D(n894), .E(n1057), .CK(clk), .Q(\mem[110][3] )
         );
  EDFFX1 \mem_reg[110][2]  ( .D(n888), .E(n1057), .CK(clk), .Q(\mem[110][2] )
         );
  EDFFX1 \mem_reg[110][1]  ( .D(n882), .E(n1057), .CK(clk), .Q(\mem[110][1] )
         );
  EDFFX1 \mem_reg[110][0]  ( .D(n876), .E(n1057), .CK(clk), .Q(\mem[110][0] )
         );
  EDFFX1 \mem_reg[114][7]  ( .D(n916), .E(n1029), .CK(clk), .Q(\mem[114][7] )
         );
  EDFFX1 \mem_reg[114][6]  ( .D(n910), .E(n1029), .CK(clk), .Q(\mem[114][6] )
         );
  EDFFX1 \mem_reg[114][5]  ( .D(n904), .E(n1029), .CK(clk), .Q(\mem[114][5] )
         );
  EDFFX1 \mem_reg[114][4]  ( .D(n898), .E(n1029), .CK(clk), .Q(\mem[114][4] )
         );
  EDFFX1 \mem_reg[114][3]  ( .D(n892), .E(n1029), .CK(clk), .Q(\mem[114][3] )
         );
  EDFFX1 \mem_reg[114][2]  ( .D(n886), .E(n1029), .CK(clk), .Q(\mem[114][2] )
         );
  EDFFX1 \mem_reg[114][1]  ( .D(n880), .E(n1029), .CK(clk), .Q(\mem[114][1] )
         );
  EDFFX1 \mem_reg[114][0]  ( .D(n874), .E(n1029), .CK(clk), .Q(\mem[114][0] )
         );
  EDFFX1 \mem_reg[118][7]  ( .D(n917), .E(n1038), .CK(clk), .Q(\mem[118][7] )
         );
  EDFFX1 \mem_reg[118][6]  ( .D(n911), .E(n1038), .CK(clk), .Q(\mem[118][6] )
         );
  EDFFX1 \mem_reg[118][5]  ( .D(n905), .E(n1038), .CK(clk), .Q(\mem[118][5] )
         );
  EDFFX1 \mem_reg[118][4]  ( .D(n899), .E(n1038), .CK(clk), .Q(\mem[118][4] )
         );
  EDFFX1 \mem_reg[118][3]  ( .D(n893), .E(n1038), .CK(clk), .Q(\mem[118][3] )
         );
  EDFFX1 \mem_reg[118][2]  ( .D(n887), .E(n1038), .CK(clk), .Q(\mem[118][2] )
         );
  EDFFX1 \mem_reg[118][1]  ( .D(n881), .E(n1038), .CK(clk), .Q(\mem[118][1] )
         );
  EDFFX1 \mem_reg[118][0]  ( .D(n875), .E(n1038), .CK(clk), .Q(\mem[118][0] )
         );
  EDFFX1 \mem_reg[122][7]  ( .D(n918), .E(n1047), .CK(clk), .Q(\mem[122][7] )
         );
  EDFFX1 \mem_reg[122][6]  ( .D(n912), .E(n1047), .CK(clk), .Q(\mem[122][6] )
         );
  EDFFX1 \mem_reg[122][5]  ( .D(n906), .E(n1047), .CK(clk), .Q(\mem[122][5] )
         );
  EDFFX1 \mem_reg[122][4]  ( .D(n900), .E(n1047), .CK(clk), .Q(\mem[122][4] )
         );
  EDFFX1 \mem_reg[122][3]  ( .D(n894), .E(n1047), .CK(clk), .Q(\mem[122][3] )
         );
  EDFFX1 \mem_reg[122][2]  ( .D(n888), .E(n1047), .CK(clk), .Q(\mem[122][2] )
         );
  EDFFX1 \mem_reg[122][1]  ( .D(n882), .E(n1047), .CK(clk), .Q(\mem[122][1] )
         );
  EDFFX1 \mem_reg[122][0]  ( .D(n876), .E(n1047), .CK(clk), .Q(\mem[122][0] )
         );
  EDFFX1 \mem_reg[126][7]  ( .D(n916), .E(n1056), .CK(clk), .Q(\mem[126][7] )
         );
  EDFFX1 \mem_reg[126][6]  ( .D(n910), .E(n1056), .CK(clk), .Q(\mem[126][6] )
         );
  EDFFX1 \mem_reg[126][5]  ( .D(n904), .E(n1056), .CK(clk), .Q(\mem[126][5] )
         );
  EDFFX1 \mem_reg[126][4]  ( .D(n898), .E(n1056), .CK(clk), .Q(\mem[126][4] )
         );
  EDFFX1 \mem_reg[126][3]  ( .D(n892), .E(n1056), .CK(clk), .Q(\mem[126][3] )
         );
  EDFFX1 \mem_reg[126][2]  ( .D(n886), .E(n1056), .CK(clk), .Q(\mem[126][2] )
         );
  EDFFX1 \mem_reg[126][1]  ( .D(n880), .E(n1056), .CK(clk), .Q(\mem[126][1] )
         );
  EDFFX1 \mem_reg[126][0]  ( .D(n874), .E(n1056), .CK(clk), .Q(\mem[126][0] )
         );
  DFFRX1 \valid_mem_reg[48]  ( .D(n1118), .CK(clk), .RN(n3), .Q(valid_mem[48])
         );
  DFFRX1 \valid_mem_reg[112]  ( .D(n1182), .CK(clk), .RN(n4), .Q(
        valid_mem[112]) );
  DFFRX1 \valid_mem_reg[49]  ( .D(n1119), .CK(clk), .RN(n3), .Q(valid_mem[49])
         );
  DFFRX1 \valid_mem_reg[113]  ( .D(n1183), .CK(clk), .RN(n4), .Q(
        valid_mem[113]) );
  DFFRX1 \valid_mem_reg[50]  ( .D(n1120), .CK(clk), .RN(n3), .Q(valid_mem[50])
         );
  DFFRX1 \valid_mem_reg[61]  ( .D(n1131), .CK(clk), .RN(n4), .Q(valid_mem[61])
         );
  DFFRX1 \valid_mem_reg[60]  ( .D(n1130), .CK(clk), .RN(n3), .Q(valid_mem[60])
         );
  DFFRX1 \valid_mem_reg[51]  ( .D(n1121), .CK(clk), .RN(n4), .Q(valid_mem[51])
         );
  DFFRX1 \valid_mem_reg[114]  ( .D(n1184), .CK(clk), .RN(n3), .Q(
        valid_mem[114]) );
  DFFRX1 \valid_mem_reg[125]  ( .D(n1195), .CK(clk), .RN(n4), .Q(
        valid_mem[125]) );
  DFFRX1 \valid_mem_reg[124]  ( .D(n1194), .CK(clk), .RN(n3), .Q(
        valid_mem[124]) );
  DFFRX1 \valid_mem_reg[115]  ( .D(n1185), .CK(clk), .RN(n4), .Q(
        valid_mem[115]) );
  DFFRX1 \valid_mem_reg[59]  ( .D(n1129), .CK(clk), .RN(n3), .Q(valid_mem[59])
         );
  DFFRX1 \valid_mem_reg[58]  ( .D(n1128), .CK(clk), .RN(n4), .Q(valid_mem[58])
         );
  DFFRX1 \valid_mem_reg[57]  ( .D(n1127), .CK(clk), .RN(n3), .Q(valid_mem[57])
         );
  DFFRX1 \valid_mem_reg[56]  ( .D(n1126), .CK(clk), .RN(n4), .Q(valid_mem[56])
         );
  DFFRX1 \valid_mem_reg[55]  ( .D(n1125), .CK(clk), .RN(n3), .Q(valid_mem[55])
         );
  DFFRX1 \valid_mem_reg[54]  ( .D(n1124), .CK(clk), .RN(n4), .Q(valid_mem[54])
         );
  DFFRX1 \valid_mem_reg[53]  ( .D(n1123), .CK(clk), .RN(n3), .Q(valid_mem[53])
         );
  DFFRX1 \valid_mem_reg[52]  ( .D(n1122), .CK(clk), .RN(n4), .Q(valid_mem[52])
         );
  DFFRX1 \valid_mem_reg[123]  ( .D(n1193), .CK(clk), .RN(n3), .Q(
        valid_mem[123]) );
  DFFRX1 \valid_mem_reg[122]  ( .D(n1192), .CK(clk), .RN(n4), .Q(
        valid_mem[122]) );
  DFFRX1 \valid_mem_reg[121]  ( .D(n1191), .CK(clk), .RN(n3), .Q(
        valid_mem[121]) );
  DFFRX1 \valid_mem_reg[120]  ( .D(n1190), .CK(clk), .RN(n4), .Q(
        valid_mem[120]) );
  DFFRX1 \valid_mem_reg[119]  ( .D(n1189), .CK(clk), .RN(n3), .Q(
        valid_mem[119]) );
  DFFRX1 \valid_mem_reg[118]  ( .D(n1188), .CK(clk), .RN(n4), .Q(
        valid_mem[118]) );
  DFFRX1 \valid_mem_reg[117]  ( .D(n1187), .CK(clk), .RN(n3), .Q(
        valid_mem[117]) );
  DFFRX1 \valid_mem_reg[116]  ( .D(n1186), .CK(clk), .RN(n4), .Q(
        valid_mem[116]) );
  DFFRX1 \valid_mem_reg[127]  ( .D(n1197), .CK(clk), .RN(n3), .Q(
        valid_mem[127]) );
  DFFRX1 \valid_mem_reg[63]  ( .D(n1133), .CK(clk), .RN(n4), .Q(valid_mem[63])
         );
  DFFRX1 \valid_mem_reg[62]  ( .D(n1132), .CK(clk), .RN(n3), .Q(valid_mem[62])
         );
  DFFRX1 \valid_mem_reg[126]  ( .D(n1196), .CK(clk), .RN(n4), .Q(
        valid_mem[126]) );
  DFFRX1 \valid_mem_reg[95]  ( .D(n1165), .CK(clk), .RN(n3), .Q(valid_mem[95])
         );
  DFFRX1 \valid_mem_reg[94]  ( .D(n1164), .CK(clk), .RN(n4), .Q(valid_mem[94])
         );
  DFFRX1 \valid_mem_reg[93]  ( .D(n1163), .CK(clk), .RN(n3), .Q(valid_mem[93])
         );
  DFFRX1 \valid_mem_reg[92]  ( .D(n1162), .CK(clk), .RN(n4), .Q(valid_mem[92])
         );
  DFFRX1 \valid_mem_reg[91]  ( .D(n1161), .CK(clk), .RN(n3), .Q(valid_mem[91])
         );
  DFFRX1 \valid_mem_reg[90]  ( .D(n1160), .CK(clk), .RN(n4), .Q(valid_mem[90])
         );
  DFFRX1 \valid_mem_reg[89]  ( .D(n1159), .CK(clk), .RN(n3), .Q(valid_mem[89])
         );
  DFFRX1 \valid_mem_reg[88]  ( .D(n1158), .CK(clk), .RN(n4), .Q(valid_mem[88])
         );
  DFFRX1 \valid_mem_reg[87]  ( .D(n1157), .CK(clk), .RN(n3), .Q(valid_mem[87])
         );
  DFFRX1 \valid_mem_reg[86]  ( .D(n1156), .CK(clk), .RN(n4), .Q(valid_mem[86])
         );
  DFFRX1 \valid_mem_reg[85]  ( .D(n1155), .CK(clk), .RN(n3), .Q(valid_mem[85])
         );
  DFFRX1 \valid_mem_reg[84]  ( .D(n1154), .CK(clk), .RN(n4), .Q(valid_mem[84])
         );
  DFFRX1 \valid_mem_reg[83]  ( .D(n1153), .CK(clk), .RN(n3), .Q(valid_mem[83])
         );
  DFFRX1 \valid_mem_reg[82]  ( .D(n1152), .CK(clk), .RN(n4), .Q(valid_mem[82])
         );
  DFFRX1 \valid_mem_reg[81]  ( .D(n1151), .CK(clk), .RN(n3), .Q(valid_mem[81])
         );
  DFFRX1 \valid_mem_reg[80]  ( .D(n1150), .CK(clk), .RN(n4), .Q(valid_mem[80])
         );
  DFFRX1 \valid_mem_reg[79]  ( .D(n1149), .CK(clk), .RN(n3), .Q(valid_mem[79])
         );
  DFFRX1 \valid_mem_reg[78]  ( .D(n1148), .CK(clk), .RN(n4), .Q(valid_mem[78])
         );
  DFFRX1 \valid_mem_reg[77]  ( .D(n1147), .CK(clk), .RN(n3), .Q(valid_mem[77])
         );
  DFFRX1 \valid_mem_reg[76]  ( .D(n1146), .CK(clk), .RN(n4), .Q(valid_mem[76])
         );
  DFFRX1 \valid_mem_reg[75]  ( .D(n1145), .CK(clk), .RN(n3), .Q(valid_mem[75])
         );
  DFFRX1 \valid_mem_reg[74]  ( .D(n1144), .CK(clk), .RN(n4), .Q(valid_mem[74])
         );
  DFFRX1 \valid_mem_reg[73]  ( .D(n1143), .CK(clk), .RN(n3), .Q(valid_mem[73])
         );
  DFFRX1 \valid_mem_reg[72]  ( .D(n1142), .CK(clk), .RN(n4), .Q(valid_mem[72])
         );
  DFFRX1 \valid_mem_reg[71]  ( .D(n1141), .CK(clk), .RN(n3), .Q(valid_mem[71])
         );
  DFFRX1 \valid_mem_reg[70]  ( .D(n1140), .CK(clk), .RN(n4), .Q(valid_mem[70])
         );
  DFFRX1 \valid_mem_reg[69]  ( .D(n1139), .CK(clk), .RN(n3), .Q(valid_mem[69])
         );
  DFFRX1 \valid_mem_reg[68]  ( .D(n1138), .CK(clk), .RN(n4), .Q(valid_mem[68])
         );
  DFFRX1 \valid_mem_reg[67]  ( .D(n1137), .CK(clk), .RN(n3), .Q(valid_mem[67])
         );
  DFFRX1 \valid_mem_reg[66]  ( .D(n1136), .CK(clk), .RN(n4), .Q(valid_mem[66])
         );
  DFFRX1 \valid_mem_reg[65]  ( .D(n1135), .CK(clk), .RN(n3), .Q(valid_mem[65])
         );
  DFFRX1 \valid_mem_reg[64]  ( .D(n1134), .CK(clk), .RN(n4), .Q(valid_mem[64])
         );
  DFFRX1 \valid_mem_reg[111]  ( .D(n1181), .CK(clk), .RN(n3), .Q(
        valid_mem[111]) );
  DFFRX1 \valid_mem_reg[110]  ( .D(n1180), .CK(clk), .RN(n4), .Q(
        valid_mem[110]) );
  DFFRX1 \valid_mem_reg[109]  ( .D(n1179), .CK(clk), .RN(n3), .Q(
        valid_mem[109]) );
  DFFRX1 \valid_mem_reg[108]  ( .D(n1178), .CK(clk), .RN(n4), .Q(
        valid_mem[108]) );
  DFFRX1 \valid_mem_reg[107]  ( .D(n1177), .CK(clk), .RN(n3), .Q(
        valid_mem[107]) );
  DFFRX1 \valid_mem_reg[106]  ( .D(n1176), .CK(clk), .RN(n4), .Q(
        valid_mem[106]) );
  DFFRX1 \valid_mem_reg[105]  ( .D(n1175), .CK(clk), .RN(n3), .Q(
        valid_mem[105]) );
  DFFRX1 \valid_mem_reg[104]  ( .D(n1174), .CK(clk), .RN(n4), .Q(
        valid_mem[104]) );
  DFFRX1 \valid_mem_reg[103]  ( .D(n1173), .CK(clk), .RN(n3), .Q(
        valid_mem[103]) );
  DFFRX1 \valid_mem_reg[102]  ( .D(n1172), .CK(clk), .RN(n4), .Q(
        valid_mem[102]) );
  DFFRX1 \valid_mem_reg[101]  ( .D(n1171), .CK(clk), .RN(n3), .Q(
        valid_mem[101]) );
  DFFRX1 \valid_mem_reg[100]  ( .D(n1170), .CK(clk), .RN(n4), .Q(
        valid_mem[100]) );
  DFFRX1 \valid_mem_reg[99]  ( .D(n1169), .CK(clk), .RN(n3), .Q(valid_mem[99])
         );
  DFFRX1 \valid_mem_reg[98]  ( .D(n1168), .CK(clk), .RN(n4), .Q(valid_mem[98])
         );
  DFFRX1 \valid_mem_reg[97]  ( .D(n1167), .CK(clk), .RN(n3), .Q(valid_mem[97])
         );
  DFFRX1 \valid_mem_reg[96]  ( .D(n1166), .CK(clk), .RN(n4), .Q(valid_mem[96])
         );
  DFFRX1 \valid_mem_reg[31]  ( .D(n1101), .CK(clk), .RN(n3), .Q(valid_mem[31])
         );
  DFFRX1 \valid_mem_reg[30]  ( .D(n1100), .CK(clk), .RN(n4), .Q(valid_mem[30])
         );
  DFFRX1 \valid_mem_reg[29]  ( .D(n1099), .CK(clk), .RN(n3), .Q(valid_mem[29])
         );
  DFFRX1 \valid_mem_reg[28]  ( .D(n1098), .CK(clk), .RN(n4), .Q(valid_mem[28])
         );
  DFFRX1 \valid_mem_reg[27]  ( .D(n1097), .CK(clk), .RN(n3), .Q(valid_mem[27])
         );
  DFFRX1 \valid_mem_reg[26]  ( .D(n1096), .CK(clk), .RN(n4), .Q(valid_mem[26])
         );
  DFFRX1 \valid_mem_reg[25]  ( .D(n1095), .CK(clk), .RN(n3), .Q(valid_mem[25])
         );
  DFFRX1 \valid_mem_reg[24]  ( .D(n1094), .CK(clk), .RN(n4), .Q(valid_mem[24])
         );
  DFFRX1 \valid_mem_reg[23]  ( .D(n1093), .CK(clk), .RN(n3), .Q(valid_mem[23])
         );
  DFFRX1 \valid_mem_reg[22]  ( .D(n1092), .CK(clk), .RN(n4), .Q(valid_mem[22])
         );
  DFFRX1 \valid_mem_reg[21]  ( .D(n1091), .CK(clk), .RN(n3), .Q(valid_mem[21])
         );
  DFFRX1 \valid_mem_reg[20]  ( .D(n1090), .CK(clk), .RN(n4), .Q(valid_mem[20])
         );
  DFFRX1 \valid_mem_reg[19]  ( .D(n1089), .CK(clk), .RN(n3), .Q(valid_mem[19])
         );
  DFFRX1 \valid_mem_reg[18]  ( .D(n1088), .CK(clk), .RN(n4), .Q(valid_mem[18])
         );
  DFFRX1 \valid_mem_reg[17]  ( .D(n1087), .CK(clk), .RN(n3), .Q(valid_mem[17])
         );
  DFFRX1 \valid_mem_reg[16]  ( .D(n1086), .CK(clk), .RN(n4), .Q(valid_mem[16])
         );
  DFFRX1 \valid_mem_reg[47]  ( .D(n1117), .CK(clk), .RN(n3), .Q(valid_mem[47])
         );
  DFFRX1 \valid_mem_reg[46]  ( .D(n1116), .CK(clk), .RN(n4), .Q(valid_mem[46])
         );
  DFFRX1 \valid_mem_reg[45]  ( .D(n1115), .CK(clk), .RN(n3), .Q(valid_mem[45])
         );
  DFFRX1 \valid_mem_reg[44]  ( .D(n1114), .CK(clk), .RN(n4), .Q(valid_mem[44])
         );
  DFFRX1 \valid_mem_reg[43]  ( .D(n1113), .CK(clk), .RN(n3), .Q(valid_mem[43])
         );
  DFFRX1 \valid_mem_reg[42]  ( .D(n1112), .CK(clk), .RN(n4), .Q(valid_mem[42])
         );
  DFFRX1 \valid_mem_reg[41]  ( .D(n1111), .CK(clk), .RN(n3), .Q(valid_mem[41])
         );
  DFFRX1 \valid_mem_reg[40]  ( .D(n1110), .CK(clk), .RN(n4), .Q(valid_mem[40])
         );
  DFFRX1 \valid_mem_reg[39]  ( .D(n1109), .CK(clk), .RN(n3), .Q(valid_mem[39])
         );
  DFFRX1 \valid_mem_reg[38]  ( .D(n1108), .CK(clk), .RN(n4), .Q(valid_mem[38])
         );
  DFFRX1 \valid_mem_reg[37]  ( .D(n1107), .CK(clk), .RN(n3), .Q(valid_mem[37])
         );
  DFFRX1 \valid_mem_reg[36]  ( .D(n1106), .CK(clk), .RN(n4), .Q(valid_mem[36])
         );
  DFFRX1 \valid_mem_reg[35]  ( .D(n1105), .CK(clk), .RN(n3), .Q(valid_mem[35])
         );
  DFFRX1 \valid_mem_reg[34]  ( .D(n1104), .CK(clk), .RN(n4), .Q(valid_mem[34])
         );
  DFFRX1 \valid_mem_reg[33]  ( .D(n1103), .CK(clk), .RN(n3), .Q(valid_mem[33])
         );
  DFFRX1 \valid_mem_reg[32]  ( .D(n1102), .CK(clk), .RN(n4), .Q(valid_mem[32])
         );
  DFFRX1 \valid_mem_reg[15]  ( .D(n1085), .CK(clk), .RN(n3), .Q(valid_mem[15])
         );
  DFFRX1 \valid_mem_reg[14]  ( .D(n1084), .CK(clk), .RN(n4), .Q(valid_mem[14])
         );
  DFFRX1 \valid_mem_reg[13]  ( .D(n1083), .CK(clk), .RN(n3), .Q(valid_mem[13])
         );
  DFFRX1 \valid_mem_reg[12]  ( .D(n1082), .CK(clk), .RN(n4), .Q(valid_mem[12])
         );
  DFFRX1 \valid_mem_reg[11]  ( .D(n1081), .CK(clk), .RN(n3), .Q(valid_mem[11])
         );
  DFFRX1 \valid_mem_reg[10]  ( .D(n1080), .CK(clk), .RN(n4), .Q(valid_mem[10])
         );
  DFFRX1 \valid_mem_reg[9]  ( .D(n1079), .CK(clk), .RN(n3), .Q(valid_mem[9])
         );
  DFFRX1 \valid_mem_reg[8]  ( .D(n1078), .CK(clk), .RN(n4), .Q(valid_mem[8])
         );
  DFFRX1 \valid_mem_reg[7]  ( .D(n1077), .CK(clk), .RN(n3), .Q(valid_mem[7])
         );
  DFFRX1 \valid_mem_reg[6]  ( .D(n1076), .CK(clk), .RN(n4), .Q(valid_mem[6])
         );
  DFFRX1 \valid_mem_reg[5]  ( .D(n1075), .CK(clk), .RN(n3), .Q(valid_mem[5])
         );
  DFFRX1 \valid_mem_reg[4]  ( .D(n1074), .CK(clk), .RN(n4), .Q(valid_mem[4])
         );
  DFFRX1 \valid_mem_reg[3]  ( .D(n1073), .CK(clk), .RN(n3), .Q(valid_mem[3])
         );
  DFFRX1 \valid_mem_reg[2]  ( .D(n1072), .CK(clk), .RN(n4), .Q(valid_mem[2])
         );
  DFFRX1 \valid_mem_reg[1]  ( .D(n1071), .CK(clk), .RN(n3), .Q(valid_mem[1])
         );
  DFFRX1 \valid_mem_reg[0]  ( .D(n1070), .CK(clk), .RN(n4), .Q(valid_mem[0])
         );
  DFFRX1 valid_reg ( .D(N41), .CK(clk), .RN(n3), .QN(n1) );
  DFFRX1 \data_out_reg[7]  ( .D(N33), .CK(clk), .RN(n4), .Q(data_out[7]) );
  DFFRX1 \data_out_reg[6]  ( .D(N34), .CK(clk), .RN(n3), .Q(data_out[6]) );
  DFFRX1 \data_out_reg[5]  ( .D(N35), .CK(clk), .RN(n4), .Q(data_out[5]) );
  DFFRX1 \data_out_reg[4]  ( .D(N36), .CK(clk), .RN(n3), .Q(data_out[4]) );
  DFFRX1 \data_out_reg[3]  ( .D(N37), .CK(clk), .RN(n4), .Q(data_out[3]) );
  DFFRX1 \data_out_reg[2]  ( .D(N38), .CK(clk), .RN(n3), .Q(data_out[2]) );
  DFFRX1 \data_out_reg[1]  ( .D(N39), .CK(clk), .RN(n4), .Q(data_out[1]) );
  DFFRX1 \data_out_reg[0]  ( .D(N40), .CK(clk), .RN(n3), .Q(data_out[0]) );
  NOR2BX4 U3 ( .AN(n871), .B(n1371), .Y(n864) );
  NOR2BX4 U4 ( .AN(n871), .B(n1338), .Y(n862) );
  NOR2BX4 U5 ( .AN(n871), .B(n1305), .Y(n860) );
  NOR2BX4 U6 ( .AN(n871), .B(n1272), .Y(n858) );
  NOR2BX4 U7 ( .AN(n871), .B(n1239), .Y(n856) );
  NAND3BXL U8 ( .AN(write_counter_count[6]), .B(n1068), .C(
        write_counter_count[5]), .Y(n1305) );
  NAND3BXL U9 ( .AN(write_counter_count[6]), .B(write_counter_count[4]), .C(
        write_counter_count[5]), .Y(n1338) );
  NAND3XL U10 ( .A(write_counter_count[5]), .B(write_counter_count[4]), .C(
        write_counter_count[6]), .Y(n1486) );
  INVX1 U11 ( .A(write_counter_count[5]), .Y(n1069) );
  INVX4 U12 ( .A(n1), .Y(valid) );
  INVX12 U13 ( .A(rst), .Y(n3) );
  INVX12 U14 ( .A(rst), .Y(n4) );
  NOR2X1 U15 ( .A(n1065), .B(n992), .Y(n1204) );
  NOR2X1 U16 ( .A(n1067), .B(n1066), .Y(n1205) );
  CLKBUFX3 U17 ( .A(n1207), .Y(n868) );
  CLKBUFX3 U18 ( .A(n1206), .Y(n866) );
  CLKBUFX3 U19 ( .A(n1208), .Y(n870) );
  NOR2X1 U20 ( .A(n1065), .B(write_counter_count[0]), .Y(n1203) );
  NOR2X1 U21 ( .A(n1066), .B(write_counter_count[3]), .Y(n1199) );
  NOR2X1 U22 ( .A(n1067), .B(write_counter_count[2]), .Y(n1200) );
  NOR2X1 U23 ( .A(n992), .B(write_counter_count[1]), .Y(n1202) );
  NOR2X1 U24 ( .A(write_counter_count[0]), .B(write_counter_count[1]), .Y(
        n1201) );
  NOR2X1 U25 ( .A(write_counter_count[2]), .B(write_counter_count[3]), .Y(
        n1198) );
  CLKBUFX3 U26 ( .A(n826), .Y(n841) );
  CLKBUFX3 U27 ( .A(n828), .Y(n838) );
  CLKBUFX3 U28 ( .A(n827), .Y(n840) );
  CLKBUFX3 U29 ( .A(n828), .Y(n839) );
  CLKBUFX3 U30 ( .A(n828), .Y(n836) );
  CLKBUFX3 U31 ( .A(n828), .Y(n837) );
  CLKBUFX3 U32 ( .A(n829), .Y(n835) );
  CLKBUFX3 U33 ( .A(n829), .Y(n834) );
  CLKBUFX3 U34 ( .A(n826), .Y(n833) );
  CLKBUFX3 U35 ( .A(n829), .Y(n831) );
  CLKBUFX3 U36 ( .A(n829), .Y(n832) );
  CLKBUFX3 U37 ( .A(n829), .Y(n830) );
  CLKBUFX3 U38 ( .A(n803), .Y(n823) );
  CLKBUFX3 U39 ( .A(n804), .Y(n821) );
  CLKBUFX3 U40 ( .A(n803), .Y(n822) );
  CLKBUFX3 U41 ( .A(n803), .Y(n818) );
  CLKBUFX3 U42 ( .A(n804), .Y(n820) );
  CLKBUFX3 U43 ( .A(n803), .Y(n819) );
  CLKBUFX3 U44 ( .A(n803), .Y(n816) );
  CLKBUFX3 U45 ( .A(n803), .Y(n817) );
  CLKBUFX3 U46 ( .A(n803), .Y(n815) );
  CLKBUFX3 U47 ( .A(n802), .Y(n814) );
  CLKBUFX3 U48 ( .A(n803), .Y(n811) );
  CLKBUFX3 U49 ( .A(n805), .Y(n813) );
  CLKBUFX3 U50 ( .A(n804), .Y(n812) );
  CLKBUFX3 U51 ( .A(n804), .Y(n809) );
  CLKBUFX3 U52 ( .A(n804), .Y(n810) );
  CLKBUFX3 U53 ( .A(n805), .Y(n806) );
  CLKBUFX3 U54 ( .A(n803), .Y(n807) );
  CLKBUFX3 U55 ( .A(n804), .Y(n808) );
  CLKBUFX3 U56 ( .A(n827), .Y(n842) );
  CLKBUFX3 U57 ( .A(n825), .Y(n827) );
  CLKBUFX3 U58 ( .A(n825), .Y(n828) );
  CLKBUFX3 U59 ( .A(n825), .Y(n829) );
  INVX3 U60 ( .A(n1485), .Y(n955) );
  INVX3 U61 ( .A(n1488), .Y(n947) );
  INVX3 U62 ( .A(n1439), .Y(n948) );
  INVX3 U63 ( .A(n1436), .Y(n1057) );
  INVX3 U64 ( .A(n1434), .Y(n984) );
  INVX3 U65 ( .A(n1432), .Y(n1021) );
  INVX3 U66 ( .A(n1430), .Y(n939) );
  INVX3 U67 ( .A(n1428), .Y(n1048) );
  INVX3 U68 ( .A(n1426), .Y(n975) );
  INVX3 U69 ( .A(n1424), .Y(n1012) );
  INVX3 U70 ( .A(n1422), .Y(n930) );
  INVX3 U71 ( .A(n1420), .Y(n1039) );
  INVX3 U72 ( .A(n1418), .Y(n966) );
  INVX3 U73 ( .A(n1416), .Y(n1003) );
  INVX3 U74 ( .A(n1414), .Y(n921) );
  INVX3 U75 ( .A(n1412), .Y(n1030) );
  INVX3 U76 ( .A(n1410), .Y(n957) );
  INVX3 U77 ( .A(n1408), .Y(n994) );
  INVX3 U78 ( .A(n1406), .Y(n949) );
  INVX3 U79 ( .A(n1403), .Y(n1058) );
  INVX3 U80 ( .A(n1401), .Y(n985) );
  INVX3 U81 ( .A(n1399), .Y(n1022) );
  INVX3 U82 ( .A(n1397), .Y(n940) );
  INVX3 U83 ( .A(n1395), .Y(n1049) );
  INVX3 U84 ( .A(n1393), .Y(n976) );
  INVX3 U85 ( .A(n1391), .Y(n1013) );
  INVX3 U86 ( .A(n1389), .Y(n931) );
  INVX3 U87 ( .A(n1387), .Y(n1040) );
  INVX3 U88 ( .A(n1385), .Y(n967) );
  INVX3 U89 ( .A(n1383), .Y(n1004) );
  INVX3 U90 ( .A(n1381), .Y(n922) );
  INVX3 U91 ( .A(n1379), .Y(n1031) );
  INVX3 U92 ( .A(n1377), .Y(n958) );
  INVX3 U93 ( .A(n1375), .Y(n995) );
  INVX3 U94 ( .A(n1373), .Y(n950) );
  INVX3 U95 ( .A(n1370), .Y(n1059) );
  INVX3 U96 ( .A(n1368), .Y(n986) );
  INVX3 U97 ( .A(n1366), .Y(n1023) );
  INVX3 U98 ( .A(n1364), .Y(n941) );
  INVX3 U99 ( .A(n1362), .Y(n1050) );
  INVX3 U100 ( .A(n1360), .Y(n977) );
  INVX3 U101 ( .A(n1358), .Y(n1014) );
  INVX3 U102 ( .A(n1356), .Y(n932) );
  INVX3 U103 ( .A(n1354), .Y(n1041) );
  INVX3 U104 ( .A(n1352), .Y(n968) );
  INVX3 U105 ( .A(n1350), .Y(n1005) );
  INVX3 U106 ( .A(n1348), .Y(n923) );
  INVX3 U107 ( .A(n1346), .Y(n1032) );
  INVX3 U108 ( .A(n1344), .Y(n959) );
  INVX3 U109 ( .A(n1342), .Y(n996) );
  INVX3 U110 ( .A(n1340), .Y(n951) );
  INVX3 U111 ( .A(n1337), .Y(n1060) );
  INVX3 U112 ( .A(n1335), .Y(n987) );
  INVX3 U113 ( .A(n1333), .Y(n1024) );
  INVX3 U114 ( .A(n1331), .Y(n942) );
  INVX3 U115 ( .A(n1329), .Y(n1051) );
  INVX3 U116 ( .A(n1327), .Y(n978) );
  INVX3 U117 ( .A(n1325), .Y(n1015) );
  INVX3 U118 ( .A(n1323), .Y(n933) );
  INVX3 U119 ( .A(n1321), .Y(n1042) );
  INVX3 U120 ( .A(n1319), .Y(n969) );
  INVX3 U121 ( .A(n1317), .Y(n1006) );
  INVX3 U122 ( .A(n1315), .Y(n924) );
  INVX3 U123 ( .A(n1313), .Y(n1033) );
  INVX3 U124 ( .A(n1311), .Y(n960) );
  INVX3 U125 ( .A(n1309), .Y(n997) );
  INVX3 U126 ( .A(n1307), .Y(n952) );
  INVX3 U127 ( .A(n1304), .Y(n1061) );
  INVX3 U128 ( .A(n1302), .Y(n988) );
  INVX3 U129 ( .A(n1300), .Y(n1025) );
  INVX3 U130 ( .A(n1298), .Y(n943) );
  INVX3 U131 ( .A(n1296), .Y(n1052) );
  INVX3 U132 ( .A(n1294), .Y(n979) );
  INVX3 U133 ( .A(n1292), .Y(n1016) );
  INVX3 U134 ( .A(n1290), .Y(n934) );
  INVX3 U135 ( .A(n1288), .Y(n1043) );
  INVX3 U136 ( .A(n1286), .Y(n970) );
  INVX3 U137 ( .A(n1284), .Y(n1007) );
  INVX3 U138 ( .A(n1282), .Y(n925) );
  INVX3 U139 ( .A(n1280), .Y(n1034) );
  INVX3 U140 ( .A(n1278), .Y(n961) );
  INVX3 U141 ( .A(n1276), .Y(n998) );
  INVX3 U142 ( .A(n1274), .Y(n953) );
  INVX3 U143 ( .A(n1271), .Y(n1062) );
  INVX3 U144 ( .A(n1269), .Y(n989) );
  INVX3 U145 ( .A(n1267), .Y(n1026) );
  INVX3 U146 ( .A(n1265), .Y(n944) );
  INVX3 U147 ( .A(n1263), .Y(n1053) );
  INVX3 U148 ( .A(n1261), .Y(n980) );
  INVX3 U149 ( .A(n1259), .Y(n1017) );
  INVX3 U150 ( .A(n1257), .Y(n935) );
  INVX3 U151 ( .A(n1255), .Y(n1044) );
  INVX3 U152 ( .A(n1253), .Y(n971) );
  INVX3 U153 ( .A(n1251), .Y(n1008) );
  INVX3 U154 ( .A(n1249), .Y(n926) );
  INVX3 U155 ( .A(n1247), .Y(n1035) );
  INVX3 U156 ( .A(n1245), .Y(n962) );
  INVX3 U157 ( .A(n1243), .Y(n999) );
  INVX3 U158 ( .A(n1241), .Y(n954) );
  INVX3 U159 ( .A(n1238), .Y(n1063) );
  INVX3 U160 ( .A(n1236), .Y(n990) );
  INVX3 U161 ( .A(n1234), .Y(n1027) );
  INVX3 U162 ( .A(n1232), .Y(n945) );
  INVX3 U163 ( .A(n1230), .Y(n1054) );
  INVX3 U164 ( .A(n1228), .Y(n981) );
  INVX3 U165 ( .A(n1226), .Y(n1018) );
  INVX3 U166 ( .A(n1224), .Y(n936) );
  INVX3 U167 ( .A(n1222), .Y(n1045) );
  INVX3 U168 ( .A(n1220), .Y(n972) );
  INVX3 U169 ( .A(n1218), .Y(n1009) );
  INVX3 U170 ( .A(n1216), .Y(n927) );
  INVX3 U171 ( .A(n1214), .Y(n1036) );
  INVX3 U172 ( .A(n1212), .Y(n963) );
  INVX3 U173 ( .A(n1210), .Y(n1000) );
  INVX3 U174 ( .A(n1484), .Y(n1056) );
  INVX3 U175 ( .A(n1481), .Y(n983) );
  INVX3 U176 ( .A(n1478), .Y(n1020) );
  INVX3 U177 ( .A(n1475), .Y(n938) );
  INVX3 U178 ( .A(n1472), .Y(n1047) );
  INVX3 U179 ( .A(n1469), .Y(n974) );
  INVX3 U180 ( .A(n1466), .Y(n1011) );
  INVX3 U181 ( .A(n1463), .Y(n929) );
  INVX3 U182 ( .A(n1460), .Y(n1038) );
  INVX3 U183 ( .A(n1457), .Y(n965) );
  INVX3 U184 ( .A(n1454), .Y(n1002) );
  INVX3 U185 ( .A(n1451), .Y(n920) );
  INVX3 U186 ( .A(n1448), .Y(n1029) );
  INVX3 U187 ( .A(n1445), .Y(n956) );
  INVX3 U188 ( .A(n1442), .Y(n993) );
  CLKBUFX3 U189 ( .A(n847), .Y(n851) );
  CLKBUFX3 U190 ( .A(n847), .Y(n850) );
  CLKBUFX3 U191 ( .A(n847), .Y(n849) );
  CLKBUFX3 U192 ( .A(n847), .Y(n848) );
  CLKBUFX3 U193 ( .A(n843), .Y(n846) );
  CLKBUFX3 U194 ( .A(n843), .Y(n845) );
  CLKBUFX3 U195 ( .A(n843), .Y(n844) );
  CLKBUFX3 U196 ( .A(n802), .Y(n805) );
  CLKBUFX3 U197 ( .A(N27), .Y(n826) );
  CLKBUFX3 U198 ( .A(N27), .Y(n825) );
  CLKBUFX3 U199 ( .A(n804), .Y(n824) );
  CLKBUFX3 U200 ( .A(data_in[0]), .Y(n872) );
  CLKBUFX3 U201 ( .A(data_in[1]), .Y(n878) );
  CLKBUFX3 U202 ( .A(data_in[2]), .Y(n884) );
  CLKBUFX3 U203 ( .A(data_in[3]), .Y(n890) );
  CLKBUFX3 U204 ( .A(data_in[4]), .Y(n896) );
  CLKBUFX3 U205 ( .A(data_in[5]), .Y(n902) );
  CLKBUFX3 U206 ( .A(data_in[6]), .Y(n908) );
  CLKBUFX3 U207 ( .A(data_in[7]), .Y(n914) );
  CLKBUFX3 U208 ( .A(data_in[0]), .Y(n873) );
  CLKBUFX3 U209 ( .A(data_in[1]), .Y(n879) );
  CLKBUFX3 U210 ( .A(data_in[2]), .Y(n885) );
  CLKBUFX3 U211 ( .A(data_in[3]), .Y(n891) );
  CLKBUFX3 U212 ( .A(data_in[4]), .Y(n897) );
  CLKBUFX3 U213 ( .A(data_in[5]), .Y(n903) );
  CLKBUFX3 U214 ( .A(data_in[6]), .Y(n909) );
  CLKBUFX3 U215 ( .A(data_in[7]), .Y(n915) );
  CLKBUFX3 U216 ( .A(n872), .Y(n874) );
  CLKBUFX3 U217 ( .A(n878), .Y(n880) );
  CLKBUFX3 U218 ( .A(n884), .Y(n886) );
  CLKBUFX3 U219 ( .A(n890), .Y(n892) );
  CLKBUFX3 U220 ( .A(n896), .Y(n898) );
  CLKBUFX3 U221 ( .A(n902), .Y(n904) );
  CLKBUFX3 U222 ( .A(n908), .Y(n910) );
  CLKBUFX3 U223 ( .A(n914), .Y(n916) );
  CLKBUFX3 U224 ( .A(n873), .Y(n875) );
  CLKBUFX3 U225 ( .A(n879), .Y(n881) );
  CLKBUFX3 U226 ( .A(n885), .Y(n887) );
  CLKBUFX3 U227 ( .A(n891), .Y(n893) );
  CLKBUFX3 U228 ( .A(n897), .Y(n899) );
  CLKBUFX3 U229 ( .A(n903), .Y(n905) );
  CLKBUFX3 U230 ( .A(n909), .Y(n911) );
  CLKBUFX3 U231 ( .A(n915), .Y(n917) );
  CLKBUFX3 U232 ( .A(n872), .Y(n876) );
  CLKBUFX3 U233 ( .A(n878), .Y(n882) );
  CLKBUFX3 U234 ( .A(n884), .Y(n888) );
  CLKBUFX3 U235 ( .A(n890), .Y(n894) );
  CLKBUFX3 U236 ( .A(n896), .Y(n900) );
  CLKBUFX3 U237 ( .A(n902), .Y(n906) );
  CLKBUFX3 U238 ( .A(n908), .Y(n912) );
  CLKBUFX3 U239 ( .A(n914), .Y(n918) );
  CLKBUFX3 U240 ( .A(n873), .Y(n877) );
  CLKBUFX3 U241 ( .A(n879), .Y(n883) );
  CLKBUFX3 U242 ( .A(n885), .Y(n889) );
  CLKBUFX3 U243 ( .A(n891), .Y(n895) );
  CLKBUFX3 U244 ( .A(n897), .Y(n901) );
  CLKBUFX3 U245 ( .A(n903), .Y(n907) );
  CLKBUFX3 U246 ( .A(n909), .Y(n913) );
  CLKBUFX3 U247 ( .A(n915), .Y(n919) );
  INVX3 U248 ( .A(n1470), .Y(n1055) );
  INVX3 U249 ( .A(n1482), .Y(n1064) );
  INVX3 U250 ( .A(n1479), .Y(n991) );
  INVX3 U251 ( .A(n1458), .Y(n1046) );
  INVX3 U252 ( .A(n1476), .Y(n1028) );
  INVX3 U253 ( .A(n1473), .Y(n946) );
  INVX3 U254 ( .A(n1467), .Y(n982) );
  INVX3 U255 ( .A(n1464), .Y(n1019) );
  INVX3 U256 ( .A(n1461), .Y(n937) );
  INVX3 U257 ( .A(n1455), .Y(n973) );
  INVX3 U258 ( .A(n1452), .Y(n1010) );
  INVX3 U259 ( .A(n1446), .Y(n1037) );
  INVX3 U260 ( .A(n1449), .Y(n928) );
  INVX3 U261 ( .A(n1443), .Y(n964) );
  INVX3 U262 ( .A(n1440), .Y(n1001) );
  NAND2X2 U263 ( .A(n1205), .B(n1204), .Y(n1485) );
  NAND2X1 U264 ( .A(n868), .B(n1064), .Y(n1436) );
  NAND2X1 U265 ( .A(n868), .B(n991), .Y(n1434) );
  NAND2X1 U266 ( .A(n868), .B(n1028), .Y(n1432) );
  NAND2X1 U267 ( .A(n868), .B(n946), .Y(n1430) );
  NAND2X1 U268 ( .A(n868), .B(n1055), .Y(n1428) );
  NAND2X1 U269 ( .A(n868), .B(n982), .Y(n1426) );
  NAND2X1 U270 ( .A(n868), .B(n1019), .Y(n1424) );
  NAND2X1 U271 ( .A(n868), .B(n937), .Y(n1422) );
  NAND2X1 U272 ( .A(n868), .B(n1046), .Y(n1420) );
  NAND2X1 U273 ( .A(n868), .B(n973), .Y(n1418) );
  NAND2X1 U274 ( .A(n868), .B(n1010), .Y(n1416) );
  NAND2X1 U275 ( .A(n868), .B(n928), .Y(n1414) );
  NAND2X1 U276 ( .A(n868), .B(n1037), .Y(n1412) );
  NAND2X1 U277 ( .A(n868), .B(n964), .Y(n1410) );
  NAND2X1 U278 ( .A(n868), .B(n1001), .Y(n1408) );
  NAND2X1 U279 ( .A(n866), .B(n1064), .Y(n1403) );
  NAND2X1 U280 ( .A(n866), .B(n991), .Y(n1401) );
  NAND2X1 U281 ( .A(n866), .B(n1028), .Y(n1399) );
  NAND2X1 U282 ( .A(n866), .B(n946), .Y(n1397) );
  NAND2X1 U283 ( .A(n866), .B(n1055), .Y(n1395) );
  NAND2X1 U284 ( .A(n866), .B(n982), .Y(n1393) );
  NAND2X1 U285 ( .A(n866), .B(n1019), .Y(n1391) );
  NAND2X1 U286 ( .A(n866), .B(n937), .Y(n1389) );
  NAND2X1 U287 ( .A(n866), .B(n1046), .Y(n1387) );
  NAND2X1 U288 ( .A(n866), .B(n973), .Y(n1385) );
  NAND2X1 U289 ( .A(n866), .B(n1010), .Y(n1383) );
  NAND2X1 U290 ( .A(n866), .B(n928), .Y(n1381) );
  NAND2X1 U291 ( .A(n866), .B(n1037), .Y(n1379) );
  NAND2X1 U292 ( .A(n866), .B(n964), .Y(n1377) );
  NAND2X1 U293 ( .A(n866), .B(n1001), .Y(n1375) );
  NAND2X1 U294 ( .A(n864), .B(n1064), .Y(n1370) );
  NAND2X1 U295 ( .A(n864), .B(n991), .Y(n1368) );
  NAND2X1 U296 ( .A(n864), .B(n1028), .Y(n1366) );
  NAND2X1 U297 ( .A(n864), .B(n946), .Y(n1364) );
  NAND2X1 U298 ( .A(n864), .B(n1055), .Y(n1362) );
  NAND2X1 U299 ( .A(n864), .B(n982), .Y(n1360) );
  NAND2X1 U300 ( .A(n864), .B(n1019), .Y(n1358) );
  NAND2X1 U301 ( .A(n864), .B(n937), .Y(n1356) );
  NAND2X1 U302 ( .A(n864), .B(n1046), .Y(n1354) );
  NAND2X1 U303 ( .A(n864), .B(n973), .Y(n1352) );
  NAND2X1 U304 ( .A(n864), .B(n1010), .Y(n1350) );
  NAND2X1 U305 ( .A(n864), .B(n928), .Y(n1348) );
  NAND2X1 U306 ( .A(n864), .B(n1037), .Y(n1346) );
  NAND2X1 U307 ( .A(n864), .B(n964), .Y(n1344) );
  NAND2X1 U308 ( .A(n864), .B(n1001), .Y(n1342) );
  NAND2X1 U309 ( .A(n862), .B(n1064), .Y(n1337) );
  NAND2X1 U310 ( .A(n862), .B(n991), .Y(n1335) );
  NAND2X1 U311 ( .A(n862), .B(n1028), .Y(n1333) );
  NAND2X1 U312 ( .A(n862), .B(n946), .Y(n1331) );
  NAND2X1 U313 ( .A(n862), .B(n1055), .Y(n1329) );
  NAND2X1 U314 ( .A(n862), .B(n982), .Y(n1327) );
  NAND2X1 U315 ( .A(n862), .B(n1019), .Y(n1325) );
  NAND2X1 U316 ( .A(n862), .B(n937), .Y(n1323) );
  NAND2X1 U317 ( .A(n862), .B(n1046), .Y(n1321) );
  NAND2X1 U318 ( .A(n862), .B(n973), .Y(n1319) );
  NAND2X1 U319 ( .A(n862), .B(n1010), .Y(n1317) );
  NAND2X1 U320 ( .A(n862), .B(n928), .Y(n1315) );
  NAND2X1 U321 ( .A(n862), .B(n1037), .Y(n1313) );
  NAND2X1 U322 ( .A(n862), .B(n964), .Y(n1311) );
  NAND2X1 U323 ( .A(n862), .B(n1001), .Y(n1309) );
  NAND2X1 U324 ( .A(n860), .B(n1064), .Y(n1304) );
  NAND2X1 U325 ( .A(n860), .B(n991), .Y(n1302) );
  NAND2X1 U326 ( .A(n860), .B(n1028), .Y(n1300) );
  NAND2X1 U327 ( .A(n860), .B(n946), .Y(n1298) );
  NAND2X1 U328 ( .A(n860), .B(n1055), .Y(n1296) );
  NAND2X1 U329 ( .A(n860), .B(n982), .Y(n1294) );
  NAND2X1 U330 ( .A(n860), .B(n1019), .Y(n1292) );
  NAND2X1 U331 ( .A(n860), .B(n937), .Y(n1290) );
  NAND2X1 U332 ( .A(n860), .B(n1046), .Y(n1288) );
  NAND2X1 U333 ( .A(n860), .B(n973), .Y(n1286) );
  NAND2X1 U334 ( .A(n860), .B(n1010), .Y(n1284) );
  NAND2X1 U335 ( .A(n860), .B(n928), .Y(n1282) );
  NAND2X1 U336 ( .A(n860), .B(n1037), .Y(n1280) );
  NAND2X1 U337 ( .A(n860), .B(n964), .Y(n1278) );
  NAND2X1 U338 ( .A(n860), .B(n1001), .Y(n1276) );
  NAND2X1 U339 ( .A(n858), .B(n1064), .Y(n1271) );
  NAND2X1 U340 ( .A(n858), .B(n991), .Y(n1269) );
  NAND2X1 U341 ( .A(n858), .B(n1028), .Y(n1267) );
  NAND2X1 U342 ( .A(n858), .B(n946), .Y(n1265) );
  NAND2X1 U343 ( .A(n858), .B(n1055), .Y(n1263) );
  NAND2X1 U344 ( .A(n858), .B(n982), .Y(n1261) );
  NAND2X1 U345 ( .A(n858), .B(n1019), .Y(n1259) );
  NAND2X1 U346 ( .A(n858), .B(n937), .Y(n1257) );
  NAND2X1 U347 ( .A(n858), .B(n1046), .Y(n1255) );
  NAND2X1 U348 ( .A(n858), .B(n973), .Y(n1253) );
  NAND2X1 U349 ( .A(n858), .B(n1010), .Y(n1251) );
  NAND2X1 U350 ( .A(n858), .B(n928), .Y(n1249) );
  NAND2X1 U351 ( .A(n858), .B(n1037), .Y(n1247) );
  NAND2X1 U352 ( .A(n858), .B(n964), .Y(n1245) );
  NAND2X1 U353 ( .A(n858), .B(n1001), .Y(n1243) );
  NAND2X1 U354 ( .A(n856), .B(n1064), .Y(n1238) );
  NAND2X1 U355 ( .A(n856), .B(n991), .Y(n1236) );
  NAND2X1 U356 ( .A(n856), .B(n1028), .Y(n1234) );
  NAND2X1 U357 ( .A(n856), .B(n946), .Y(n1232) );
  NAND2X1 U358 ( .A(n856), .B(n1055), .Y(n1230) );
  NAND2X1 U359 ( .A(n856), .B(n982), .Y(n1228) );
  NAND2X1 U360 ( .A(n856), .B(n1019), .Y(n1226) );
  NAND2X1 U361 ( .A(n856), .B(n937), .Y(n1224) );
  NAND2X1 U362 ( .A(n856), .B(n1046), .Y(n1222) );
  NAND2X1 U363 ( .A(n856), .B(n973), .Y(n1220) );
  NAND2X1 U364 ( .A(n856), .B(n1010), .Y(n1218) );
  NAND2X1 U365 ( .A(n856), .B(n928), .Y(n1216) );
  NAND2X1 U366 ( .A(n856), .B(n1037), .Y(n1214) );
  NAND2X1 U367 ( .A(n856), .B(n964), .Y(n1212) );
  NAND2X1 U368 ( .A(n856), .B(n1001), .Y(n1210) );
  NAND2X1 U369 ( .A(n870), .B(n955), .Y(n1488) );
  NAND2X1 U370 ( .A(n868), .B(n955), .Y(n1439) );
  NAND2X1 U371 ( .A(n866), .B(n955), .Y(n1406) );
  NAND2X1 U372 ( .A(n864), .B(n955), .Y(n1373) );
  NAND2X1 U373 ( .A(n862), .B(n955), .Y(n1340) );
  NAND2X1 U374 ( .A(n860), .B(n955), .Y(n1307) );
  NAND2X1 U375 ( .A(n858), .B(n955), .Y(n1274) );
  NAND2X1 U376 ( .A(n856), .B(n955), .Y(n1241) );
  NAND2X1 U377 ( .A(n1064), .B(n870), .Y(n1484) );
  NAND2X1 U378 ( .A(n991), .B(n870), .Y(n1481) );
  NAND2X1 U379 ( .A(n1028), .B(n870), .Y(n1478) );
  NAND2X1 U380 ( .A(n946), .B(n870), .Y(n1475) );
  NAND2X1 U381 ( .A(n1055), .B(n870), .Y(n1472) );
  NAND2X1 U382 ( .A(n982), .B(n870), .Y(n1469) );
  NAND2X1 U383 ( .A(n1019), .B(n870), .Y(n1466) );
  NAND2X1 U384 ( .A(n937), .B(n870), .Y(n1463) );
  NAND2X1 U385 ( .A(n1046), .B(n870), .Y(n1460) );
  NAND2X1 U386 ( .A(n973), .B(n870), .Y(n1457) );
  NAND2X1 U387 ( .A(n1010), .B(n870), .Y(n1454) );
  NAND2X1 U388 ( .A(n928), .B(n870), .Y(n1451) );
  NAND2X1 U389 ( .A(n1037), .B(n870), .Y(n1448) );
  NAND2X1 U390 ( .A(n964), .B(n870), .Y(n1445) );
  NAND2X1 U391 ( .A(n1001), .B(n870), .Y(n1442) );
  CLKBUFX3 U392 ( .A(N29), .Y(n847) );
  CLKBUFX3 U393 ( .A(N28), .Y(n843) );
  CLKBUFX3 U394 ( .A(N26), .Y(n804) );
  CLKBUFX3 U395 ( .A(N26), .Y(n803) );
  CLKBUFX3 U396 ( .A(N26), .Y(n802) );
  NAND2X2 U397 ( .A(n1200), .B(n1203), .Y(n1470) );
  NAND2X2 U398 ( .A(n1199), .B(n1203), .Y(n1458) );
  NAND2X2 U399 ( .A(n1198), .B(n1203), .Y(n1446) );
  NAND2X2 U400 ( .A(n1200), .B(n1201), .Y(n1464) );
  NAND2X2 U401 ( .A(n1199), .B(n1201), .Y(n1452) );
  NAND2X2 U402 ( .A(n1198), .B(n1201), .Y(n1440) );
  NAND2X2 U403 ( .A(n1200), .B(n1202), .Y(n1467) );
  NAND2X2 U404 ( .A(n1199), .B(n1202), .Y(n1455) );
  NAND2X2 U405 ( .A(n1198), .B(n1202), .Y(n1443) );
  NAND2X2 U406 ( .A(n1203), .B(n1205), .Y(n1482) );
  NAND2X2 U407 ( .A(n1202), .B(n1205), .Y(n1479) );
  NAND2X2 U408 ( .A(n1201), .B(n1205), .Y(n1476) );
  NAND2X2 U409 ( .A(n1200), .B(n1204), .Y(n1473) );
  NAND2X2 U410 ( .A(n1199), .B(n1204), .Y(n1461) );
  NAND2X2 U411 ( .A(n1198), .B(n1204), .Y(n1449) );
  BUFX4 U412 ( .A(N31), .Y(n853) );
  MXI2X1 U413 ( .A(n728), .B(n729), .S0(n854), .Y(N40) );
  MX4X1 U414 ( .A(n801), .B(n799), .C(n800), .D(n798), .S0(n853), .S1(n852), 
        .Y(n728) );
  MX4X1 U415 ( .A(n797), .B(n795), .C(n796), .D(n794), .S0(n853), .S1(n852), 
        .Y(n729) );
  MXI4X1 U416 ( .A(n727), .B(n725), .C(n726), .D(n724), .S0(n851), .S1(n846), 
        .Y(n801) );
  MXI2X1 U417 ( .A(n694), .B(n695), .S0(n854), .Y(N39) );
  MX4X1 U418 ( .A(n793), .B(n791), .C(n792), .D(n790), .S0(n853), .S1(n852), 
        .Y(n694) );
  MX4X1 U419 ( .A(n789), .B(n787), .C(n788), .D(n786), .S0(n853), .S1(n852), 
        .Y(n695) );
  MXI4X1 U420 ( .A(n693), .B(n691), .C(n692), .D(n690), .S0(n851), .S1(n846), 
        .Y(n793) );
  MXI2X1 U421 ( .A(n660), .B(n661), .S0(n854), .Y(N38) );
  MX4X1 U422 ( .A(n785), .B(n783), .C(n784), .D(n782), .S0(n853), .S1(n852), 
        .Y(n660) );
  MX4X1 U423 ( .A(n781), .B(n779), .C(n780), .D(n778), .S0(n853), .S1(n852), 
        .Y(n661) );
  MXI4X1 U424 ( .A(n659), .B(n657), .C(n658), .D(n656), .S0(n850), .S1(n846), 
        .Y(n785) );
  MXI2X1 U425 ( .A(n626), .B(n627), .S0(n854), .Y(N37) );
  MX4X1 U426 ( .A(n777), .B(n775), .C(n776), .D(n774), .S0(n853), .S1(n852), 
        .Y(n626) );
  MX4X1 U427 ( .A(n773), .B(n771), .C(n772), .D(n770), .S0(n853), .S1(n852), 
        .Y(n627) );
  MXI4X1 U428 ( .A(n625), .B(n623), .C(n624), .D(n622), .S0(n849), .S1(n845), 
        .Y(n777) );
  MXI2X1 U429 ( .A(n592), .B(n593), .S0(n854), .Y(N36) );
  MX4X1 U430 ( .A(n769), .B(n767), .C(n768), .D(n766), .S0(n853), .S1(n852), 
        .Y(n592) );
  MX4X1 U431 ( .A(n765), .B(n763), .C(n764), .D(n762), .S0(n853), .S1(n852), 
        .Y(n593) );
  MXI4X1 U432 ( .A(n591), .B(n589), .C(n590), .D(n588), .S0(n849), .S1(n845), 
        .Y(n769) );
  MXI2X1 U433 ( .A(n139), .B(n140), .S0(n854), .Y(N35) );
  MX4X1 U434 ( .A(n761), .B(n759), .C(n760), .D(n758), .S0(n853), .S1(n852), 
        .Y(n139) );
  MX4X1 U435 ( .A(n757), .B(n755), .C(n756), .D(n754), .S0(n853), .S1(n852), 
        .Y(n140) );
  MXI4X1 U436 ( .A(n138), .B(n136), .C(n137), .D(n135), .S0(n849), .S1(n844), 
        .Y(n761) );
  MXI2X1 U437 ( .A(n105), .B(n106), .S0(n854), .Y(N34) );
  MX4X1 U438 ( .A(n753), .B(n751), .C(n752), .D(n750), .S0(n853), .S1(n852), 
        .Y(n105) );
  MX4X1 U439 ( .A(n749), .B(n747), .C(n748), .D(n746), .S0(n853), .S1(n852), 
        .Y(n106) );
  MXI4X1 U440 ( .A(n104), .B(n102), .C(n103), .D(n101), .S0(n847), .S1(n844), 
        .Y(n753) );
  MXI2X1 U441 ( .A(n71), .B(n72), .S0(n854), .Y(N33) );
  MX4X1 U442 ( .A(n745), .B(n743), .C(n744), .D(n742), .S0(n853), .S1(n852), 
        .Y(n71) );
  MX4X1 U443 ( .A(n741), .B(n739), .C(n740), .D(n738), .S0(n853), .S1(n852), 
        .Y(n72) );
  MXI4X1 U444 ( .A(n70), .B(n68), .C(n69), .D(n67), .S0(n847), .S1(n846), .Y(
        n745) );
  MXI2X1 U445 ( .A(n37), .B(n38), .S0(n854), .Y(N41) );
  MX4X1 U446 ( .A(n737), .B(n735), .C(n736), .D(n734), .S0(n853), .S1(n852), 
        .Y(n37) );
  MX4X1 U447 ( .A(n733), .B(n731), .C(n732), .D(n730), .S0(n853), .S1(n852), 
        .Y(n38) );
  MXI4X1 U448 ( .A(n36), .B(n34), .C(n35), .D(n33), .S0(n848), .S1(n843), .Y(
        n737) );
  NOR2BX1 U449 ( .AN(n871), .B(n867), .Y(n1207) );
  NOR2BX1 U450 ( .AN(n871), .B(n865), .Y(n1206) );
  BUFX4 U451 ( .A(N30), .Y(n852) );
  NOR2BX1 U452 ( .AN(n871), .B(n869), .Y(n1208) );
  CLKBUFX3 U453 ( .A(en), .Y(n871) );
  CLKINVX1 U454 ( .A(write_counter_count[4]), .Y(n1068) );
  CLKINVX1 U455 ( .A(write_counter_count[0]), .Y(n992) );
  CLKBUFX3 U456 ( .A(n1305), .Y(n859) );
  CLKBUFX3 U457 ( .A(n1486), .Y(n869) );
  CLKINVX1 U458 ( .A(write_counter_count[2]), .Y(n1066) );
  CLKINVX1 U459 ( .A(write_counter_count[3]), .Y(n1067) );
  CLKINVX1 U460 ( .A(write_counter_count[1]), .Y(n1065) );
  CLKBUFX3 U461 ( .A(n1338), .Y(n861) );
  CLKBUFX3 U462 ( .A(n1437), .Y(n867) );
  NAND3X1 U463 ( .A(write_counter_count[5]), .B(n1068), .C(
        write_counter_count[6]), .Y(n1437) );
  CLKBUFX3 U464 ( .A(n1404), .Y(n865) );
  NAND3X1 U465 ( .A(write_counter_count[4]), .B(n1069), .C(
        write_counter_count[6]), .Y(n1404) );
  CLKBUFX3 U466 ( .A(n1272), .Y(n857) );
  NAND3BX1 U467 ( .AN(write_counter_count[6]), .B(n1069), .C(
        write_counter_count[4]), .Y(n1272) );
  CLKBUFX3 U468 ( .A(n1371), .Y(n863) );
  NAND3X1 U469 ( .A(n1068), .B(n1069), .C(write_counter_count[6]), .Y(n1371)
         );
  CLKBUFX3 U470 ( .A(n1239), .Y(n855) );
  NAND3BX1 U471 ( .AN(write_counter_count[6]), .B(n1069), .C(n1068), .Y(n1239)
         );
  MX4X1 U472 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .C(\mem[6][0] ), .D(
        \mem[7][0] ), .S0(n824), .S1(n842), .Y(n726) );
  MX4X1 U473 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .C(\mem[6][1] ), .D(
        \mem[7][1] ), .S0(n822), .S1(n825), .Y(n692) );
  MX4X1 U474 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .C(\mem[6][2] ), .D(
        \mem[7][2] ), .S0(n819), .S1(n839), .Y(n658) );
  MX4X1 U475 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .C(\mem[6][3] ), .D(
        \mem[7][3] ), .S0(n817), .S1(n837), .Y(n624) );
  MX4X1 U476 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .C(\mem[6][4] ), .D(
        \mem[7][4] ), .S0(n815), .S1(n835), .Y(n590) );
  MX4X1 U477 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .C(\mem[6][5] ), .D(
        \mem[7][5] ), .S0(n802), .S1(n825), .Y(n137) );
  MX4X1 U478 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .C(\mem[6][6] ), .D(
        \mem[7][6] ), .S0(n813), .S1(n840), .Y(n103) );
  MX4X1 U479 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .C(\mem[6][7] ), .D(
        \mem[7][7] ), .S0(n810), .S1(n832), .Y(n69) );
  MX4X1 U480 ( .A(valid_mem[4]), .B(valid_mem[5]), .C(valid_mem[6]), .D(
        valid_mem[7]), .S0(n808), .S1(n842), .Y(n35) );
  MX4X1 U481 ( .A(\mem[80][0] ), .B(\mem[81][0] ), .C(\mem[82][0] ), .D(
        \mem[83][0] ), .S0(n823), .S1(n827), .Y(n707) );
  MX4X1 U482 ( .A(\mem[112][0] ), .B(\mem[113][0] ), .C(\mem[114][0] ), .D(
        \mem[115][0] ), .S0(n822), .S1(n835), .Y(n699) );
  MX4X1 U483 ( .A(\mem[96][0] ), .B(\mem[97][0] ), .C(\mem[98][0] ), .D(
        \mem[99][0] ), .S0(n823), .S1(n827), .Y(n703) );
  MX4X1 U484 ( .A(\mem[64][0] ), .B(\mem[65][0] ), .C(\mem[66][0] ), .D(
        \mem[67][0] ), .S0(n823), .S1(n831), .Y(n711) );
  MX4X1 U485 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .C(\mem[18][0] ), .D(
        \mem[19][0] ), .S0(n824), .S1(n842), .Y(n723) );
  MX4X1 U486 ( .A(\mem[32][0] ), .B(\mem[33][0] ), .C(\mem[34][0] ), .D(
        \mem[35][0] ), .S0(n824), .S1(n842), .Y(n719) );
  MX4X1 U487 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .C(\mem[2][0] ), .D(
        \mem[3][0] ), .S0(n824), .S1(n842), .Y(n727) );
  MX4X1 U488 ( .A(\mem[80][1] ), .B(\mem[81][1] ), .C(\mem[82][1] ), .D(
        \mem[83][1] ), .S0(n820), .S1(n840), .Y(n673) );
  MX4X1 U489 ( .A(\mem[112][1] ), .B(\mem[113][1] ), .C(\mem[114][1] ), .D(
        \mem[115][1] ), .S0(n820), .S1(n840), .Y(n665) );
  MX4X1 U490 ( .A(\mem[96][1] ), .B(\mem[97][1] ), .C(\mem[98][1] ), .D(
        \mem[99][1] ), .S0(n820), .S1(n840), .Y(n669) );
  MX4X1 U491 ( .A(\mem[64][1] ), .B(\mem[65][1] ), .C(\mem[66][1] ), .D(
        \mem[67][1] ), .S0(n821), .S1(n841), .Y(n677) );
  MX4X1 U492 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .C(\mem[18][1] ), .D(
        \mem[19][1] ), .S0(n822), .S1(n827), .Y(n689) );
  MX4X1 U493 ( .A(\mem[48][1] ), .B(\mem[49][1] ), .C(\mem[50][1] ), .D(
        \mem[51][1] ), .S0(n821), .S1(n841), .Y(n681) );
  MX4X1 U494 ( .A(\mem[32][1] ), .B(\mem[33][1] ), .C(\mem[34][1] ), .D(
        \mem[35][1] ), .S0(n821), .S1(n841), .Y(n685) );
  MX4X1 U495 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .C(\mem[2][1] ), .D(
        \mem[3][1] ), .S0(n822), .S1(n833), .Y(n693) );
  MX4X1 U496 ( .A(\mem[80][2] ), .B(\mem[81][2] ), .C(\mem[82][2] ), .D(
        \mem[83][2] ), .S0(n818), .S1(n838), .Y(n639) );
  MX4X1 U497 ( .A(\mem[112][2] ), .B(\mem[113][2] ), .C(\mem[114][2] ), .D(
        \mem[115][2] ), .S0(n817), .S1(n837), .Y(n631) );
  MX4X1 U498 ( .A(\mem[96][2] ), .B(\mem[97][2] ), .C(\mem[98][2] ), .D(
        \mem[99][2] ), .S0(n818), .S1(n838), .Y(n635) );
  MX4X1 U499 ( .A(\mem[64][2] ), .B(\mem[65][2] ), .C(\mem[66][2] ), .D(
        \mem[67][2] ), .S0(n818), .S1(n838), .Y(n643) );
  MX4X1 U500 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .C(\mem[18][2] ), .D(
        \mem[19][2] ), .S0(n819), .S1(n839), .Y(n655) );
  MX4X1 U501 ( .A(\mem[48][2] ), .B(\mem[49][2] ), .C(\mem[50][2] ), .D(
        \mem[51][2] ), .S0(n819), .S1(n839), .Y(n647) );
  MX4X1 U502 ( .A(\mem[32][2] ), .B(\mem[33][2] ), .C(\mem[34][2] ), .D(
        \mem[35][2] ), .S0(n819), .S1(n839), .Y(n651) );
  MX4X1 U503 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .C(\mem[2][2] ), .D(
        \mem[3][2] ), .S0(n820), .S1(n840), .Y(n659) );
  MX4X1 U504 ( .A(\mem[80][3] ), .B(\mem[81][3] ), .C(\mem[82][3] ), .D(
        \mem[83][3] ), .S0(n816), .S1(n836), .Y(n605) );
  MX4X1 U505 ( .A(\mem[112][3] ), .B(\mem[113][3] ), .C(\mem[114][3] ), .D(
        \mem[115][3] ), .S0(n815), .S1(n835), .Y(n597) );
  MX4X1 U506 ( .A(\mem[96][3] ), .B(\mem[97][3] ), .C(\mem[98][3] ), .D(
        \mem[99][3] ), .S0(n815), .S1(n835), .Y(n601) );
  MX4X1 U507 ( .A(\mem[64][3] ), .B(\mem[65][3] ), .C(\mem[66][3] ), .D(
        \mem[67][3] ), .S0(n816), .S1(n836), .Y(n609) );
  MX4X1 U508 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .C(\mem[18][3] ), .D(
        \mem[19][3] ), .S0(n817), .S1(n837), .Y(n621) );
  MX4X1 U509 ( .A(\mem[48][3] ), .B(\mem[49][3] ), .C(\mem[50][3] ), .D(
        \mem[51][3] ), .S0(n816), .S1(n836), .Y(n613) );
  MX4X1 U510 ( .A(\mem[32][3] ), .B(\mem[33][3] ), .C(\mem[34][3] ), .D(
        \mem[35][3] ), .S0(n816), .S1(n836), .Y(n617) );
  MX4X1 U511 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .C(\mem[2][3] ), .D(
        \mem[3][3] ), .S0(n817), .S1(n837), .Y(n625) );
  MX4X1 U512 ( .A(\mem[80][4] ), .B(\mem[81][4] ), .C(\mem[82][4] ), .D(
        \mem[83][4] ), .S0(n805), .S1(n826), .Y(n435) );
  MX4X1 U513 ( .A(\mem[112][4] ), .B(\mem[113][4] ), .C(\mem[114][4] ), .D(
        \mem[115][4] ), .S0(n804), .S1(n827), .Y(n144) );
  MX4X1 U514 ( .A(\mem[96][4] ), .B(\mem[97][4] ), .C(\mem[98][4] ), .D(
        \mem[99][4] ), .S0(n805), .S1(n825), .Y(n148) );
  MX4X1 U515 ( .A(\mem[64][4] ), .B(\mem[65][4] ), .C(\mem[66][4] ), .D(
        \mem[67][4] ), .S0(n805), .S1(n826), .Y(n439) );
  MX4X1 U516 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .C(\mem[18][4] ), .D(
        \mem[19][4] ), .S0(n803), .S1(n834), .Y(n587) );
  MX4X1 U517 ( .A(\mem[48][4] ), .B(\mem[49][4] ), .C(\mem[50][4] ), .D(
        \mem[51][4] ), .S0(n805), .S1(n834), .Y(n579) );
  MX4X1 U518 ( .A(\mem[32][4] ), .B(\mem[33][4] ), .C(\mem[34][4] ), .D(
        \mem[35][4] ), .S0(n804), .S1(n834), .Y(n583) );
  MX4X1 U519 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .C(\mem[2][4] ), .D(
        \mem[3][4] ), .S0(n815), .S1(n835), .Y(n591) );
  MX4X1 U520 ( .A(\mem[80][5] ), .B(\mem[81][5] ), .C(\mem[82][5] ), .D(
        \mem[83][5] ), .S0(n814), .S1(n840), .Y(n118) );
  MX4X1 U521 ( .A(\mem[112][5] ), .B(\mem[113][5] ), .C(\mem[114][5] ), .D(
        \mem[115][5] ), .S0(n813), .S1(n828), .Y(n110) );
  MX4X1 U522 ( .A(\mem[96][5] ), .B(\mem[97][5] ), .C(\mem[98][5] ), .D(
        \mem[99][5] ), .S0(n813), .S1(n827), .Y(n114) );
  MX4X1 U523 ( .A(\mem[64][5] ), .B(\mem[65][5] ), .C(\mem[66][5] ), .D(
        \mem[67][5] ), .S0(n814), .S1(n825), .Y(n122) );
  MX4X1 U524 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .C(\mem[18][5] ), .D(
        \mem[19][5] ), .S0(n803), .S1(n826), .Y(n134) );
  MX4X1 U525 ( .A(\mem[48][5] ), .B(\mem[49][5] ), .C(\mem[50][5] ), .D(
        \mem[51][5] ), .S0(n814), .S1(n828), .Y(n126) );
  MX4X1 U526 ( .A(\mem[32][5] ), .B(\mem[33][5] ), .C(\mem[34][5] ), .D(
        \mem[35][5] ), .S0(n802), .S1(n826), .Y(n130) );
  MX4X1 U527 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .C(\mem[2][5] ), .D(
        \mem[3][5] ), .S0(n802), .S1(n826), .Y(n138) );
  MX4X1 U528 ( .A(\mem[80][6] ), .B(\mem[81][6] ), .C(\mem[82][6] ), .D(
        \mem[83][6] ), .S0(n811), .S1(n836), .Y(n84) );
  MX4X1 U529 ( .A(\mem[112][6] ), .B(\mem[113][6] ), .C(\mem[114][6] ), .D(
        \mem[115][6] ), .S0(n811), .S1(n832), .Y(n76) );
  MX4X1 U530 ( .A(\mem[96][6] ), .B(\mem[97][6] ), .C(\mem[98][6] ), .D(
        \mem[99][6] ), .S0(n811), .S1(n826), .Y(n80) );
  MX4X1 U531 ( .A(\mem[64][6] ), .B(\mem[65][6] ), .C(\mem[66][6] ), .D(
        \mem[67][6] ), .S0(n811), .S1(n830), .Y(n88) );
  MX4X1 U532 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .C(\mem[18][6] ), .D(
        \mem[19][6] ), .S0(n812), .S1(n833), .Y(n100) );
  MX4X1 U533 ( .A(\mem[48][6] ), .B(\mem[49][6] ), .C(\mem[50][6] ), .D(
        \mem[51][6] ), .S0(n812), .S1(n833), .Y(n92) );
  MX4X1 U534 ( .A(\mem[32][6] ), .B(\mem[33][6] ), .C(\mem[34][6] ), .D(
        \mem[35][6] ), .S0(n812), .S1(n833), .Y(n96) );
  MX4X1 U535 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .C(\mem[2][6] ), .D(
        \mem[3][6] ), .S0(n813), .S1(n825), .Y(n104) );
  MX4X1 U536 ( .A(\mem[80][7] ), .B(\mem[81][7] ), .C(\mem[82][7] ), .D(
        \mem[83][7] ), .S0(n809), .S1(n831), .Y(n50) );
  MX4X1 U537 ( .A(\mem[112][7] ), .B(\mem[113][7] ), .C(\mem[114][7] ), .D(
        \mem[115][7] ), .S0(n808), .S1(n832), .Y(n42) );
  MX4X1 U538 ( .A(\mem[96][7] ), .B(\mem[97][7] ), .C(\mem[98][7] ), .D(
        \mem[99][7] ), .S0(n808), .S1(n838), .Y(n46) );
  MX4X1 U539 ( .A(\mem[64][7] ), .B(\mem[65][7] ), .C(\mem[66][7] ), .D(
        \mem[67][7] ), .S0(n809), .S1(n831), .Y(n54) );
  MX4X1 U540 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .C(\mem[18][7] ), .D(
        \mem[19][7] ), .S0(n810), .S1(n832), .Y(n66) );
  MX4X1 U541 ( .A(\mem[48][7] ), .B(\mem[49][7] ), .C(\mem[50][7] ), .D(
        \mem[51][7] ), .S0(n809), .S1(n831), .Y(n58) );
  MX4X1 U542 ( .A(\mem[32][7] ), .B(\mem[33][7] ), .C(\mem[34][7] ), .D(
        \mem[35][7] ), .S0(n810), .S1(n832), .Y(n62) );
  MX4X1 U543 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .C(\mem[2][7] ), .D(
        \mem[3][7] ), .S0(n810), .S1(n832), .Y(n70) );
  MX4X1 U544 ( .A(valid_mem[80]), .B(valid_mem[81]), .C(valid_mem[82]), .D(
        valid_mem[83]), .S0(n806), .S1(n839), .Y(n16) );
  MX4X1 U545 ( .A(valid_mem[112]), .B(valid_mem[113]), .C(valid_mem[114]), .D(
        valid_mem[115]), .S0(n806), .S1(n840), .Y(n8) );
  MX4X1 U546 ( .A(valid_mem[96]), .B(valid_mem[97]), .C(valid_mem[98]), .D(
        valid_mem[99]), .S0(n806), .S1(n825), .Y(n12) );
  MX4X1 U547 ( .A(valid_mem[64]), .B(valid_mem[65]), .C(valid_mem[66]), .D(
        valid_mem[67]), .S0(n807), .S1(n830), .Y(n20) );
  MX4X1 U548 ( .A(valid_mem[16]), .B(valid_mem[17]), .C(valid_mem[18]), .D(
        valid_mem[19]), .S0(n807), .S1(n830), .Y(n32) );
  MX4X1 U549 ( .A(valid_mem[48]), .B(valid_mem[49]), .C(valid_mem[50]), .D(
        valid_mem[51]), .S0(n807), .S1(n830), .Y(n24) );
  MX4X1 U550 ( .A(valid_mem[32]), .B(valid_mem[33]), .C(valid_mem[34]), .D(
        valid_mem[35]), .S0(n807), .S1(n830), .Y(n28) );
  MX4X1 U551 ( .A(valid_mem[0]), .B(valid_mem[1]), .C(valid_mem[2]), .D(
        valid_mem[3]), .S0(n808), .S1(n827), .Y(n36) );
  MX4X1 U552 ( .A(\mem[56][0] ), .B(\mem[57][0] ), .C(\mem[58][0] ), .D(
        \mem[59][0] ), .S0(n823), .S1(n827), .Y(n713) );
  MX4X1 U553 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .C(\mem[10][0] ), .D(
        \mem[11][0] ), .S0(n824), .S1(n842), .Y(n725) );
  MX4X1 U554 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .C(\mem[10][1] ), .D(
        \mem[11][1] ), .S0(n822), .S1(n829), .Y(n691) );
  MX4X1 U555 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .C(\mem[10][2] ), .D(
        \mem[11][2] ), .S0(n819), .S1(n839), .Y(n657) );
  MX4X1 U556 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .C(\mem[10][3] ), .D(
        \mem[11][3] ), .S0(n817), .S1(n837), .Y(n623) );
  MX4X1 U557 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .C(\mem[10][4] ), .D(
        \mem[11][4] ), .S0(N26), .S1(n834), .Y(n589) );
  MX4X1 U558 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .C(\mem[10][5] ), .D(
        \mem[11][5] ), .S0(n804), .S1(n825), .Y(n136) );
  MX4X1 U559 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .C(\mem[10][6] ), .D(
        \mem[11][6] ), .S0(n813), .S1(n826), .Y(n102) );
  MX4X1 U560 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .C(\mem[10][7] ), .D(
        \mem[11][7] ), .S0(n810), .S1(n832), .Y(n68) );
  MX4X1 U561 ( .A(valid_mem[8]), .B(valid_mem[9]), .C(valid_mem[10]), .D(
        valid_mem[11]), .S0(n808), .S1(n837), .Y(n34) );
  MX4X1 U562 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .C(\mem[14][0] ), .D(
        \mem[15][0] ), .S0(n824), .S1(n842), .Y(n724) );
  MX4X1 U563 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .C(\mem[14][1] ), .D(
        \mem[15][1] ), .S0(n822), .S1(n827), .Y(n690) );
  MX4X1 U564 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .C(\mem[14][2] ), .D(
        \mem[15][2] ), .S0(n819), .S1(n839), .Y(n656) );
  MX4X1 U565 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .C(\mem[14][3] ), .D(
        \mem[15][3] ), .S0(n817), .S1(n837), .Y(n622) );
  MX4X1 U566 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .C(\mem[14][4] ), .D(
        \mem[15][4] ), .S0(N26), .S1(n834), .Y(n588) );
  MX4X1 U567 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .C(\mem[14][5] ), .D(
        \mem[15][5] ), .S0(n802), .S1(n826), .Y(n135) );
  MX4X1 U568 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .C(\mem[14][6] ), .D(
        \mem[15][6] ), .S0(n812), .S1(n833), .Y(n101) );
  MX4X1 U569 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .C(\mem[14][7] ), .D(
        \mem[15][7] ), .S0(n810), .S1(n832), .Y(n67) );
  MX4X1 U570 ( .A(valid_mem[12]), .B(valid_mem[13]), .C(valid_mem[14]), .D(
        valid_mem[15]), .S0(n808), .S1(n840), .Y(n33) );
  CLKBUFX3 U571 ( .A(N32), .Y(n854) );
  MXI4X1 U572 ( .A(n707), .B(n705), .C(n706), .D(n704), .S0(n851), .S1(n846), 
        .Y(n796) );
  MX4X1 U573 ( .A(\mem[92][0] ), .B(\mem[93][0] ), .C(\mem[94][0] ), .D(
        \mem[95][0] ), .S0(n823), .S1(n829), .Y(n704) );
  MX4X1 U574 ( .A(\mem[84][0] ), .B(\mem[85][0] ), .C(\mem[86][0] ), .D(
        \mem[87][0] ), .S0(n823), .S1(n828), .Y(n706) );
  MX4X1 U575 ( .A(\mem[88][0] ), .B(\mem[89][0] ), .C(\mem[90][0] ), .D(
        \mem[91][0] ), .S0(n823), .S1(n828), .Y(n705) );
  MXI4X1 U576 ( .A(n723), .B(n721), .C(n722), .D(n720), .S0(n851), .S1(n846), 
        .Y(n800) );
  MX4X1 U577 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .C(\mem[30][0] ), .D(
        \mem[31][0] ), .S0(n824), .S1(n842), .Y(n720) );
  MX4X1 U578 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .C(\mem[22][0] ), .D(
        \mem[23][0] ), .S0(n824), .S1(n842), .Y(n722) );
  MX4X1 U579 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .C(\mem[26][0] ), .D(
        \mem[27][0] ), .S0(n824), .S1(n842), .Y(n721) );
  MXI4X1 U580 ( .A(n673), .B(n671), .C(n672), .D(n670), .S0(n850), .S1(n846), 
        .Y(n788) );
  MX4X1 U581 ( .A(\mem[92][1] ), .B(\mem[93][1] ), .C(\mem[94][1] ), .D(
        \mem[95][1] ), .S0(n820), .S1(n840), .Y(n670) );
  MX4X1 U582 ( .A(\mem[84][1] ), .B(\mem[85][1] ), .C(\mem[86][1] ), .D(
        \mem[87][1] ), .S0(n820), .S1(n840), .Y(n672) );
  MX4X1 U583 ( .A(\mem[88][1] ), .B(\mem[89][1] ), .C(\mem[90][1] ), .D(
        \mem[91][1] ), .S0(n820), .S1(n840), .Y(n671) );
  MXI4X1 U584 ( .A(n689), .B(n687), .C(n688), .D(n686), .S0(n851), .S1(n846), 
        .Y(n792) );
  MX4X1 U585 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .C(\mem[30][1] ), .D(
        \mem[31][1] ), .S0(n821), .S1(n841), .Y(n686) );
  MX4X1 U586 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .C(\mem[22][1] ), .D(
        \mem[23][1] ), .S0(n822), .S1(n826), .Y(n688) );
  MX4X1 U587 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .C(\mem[26][1] ), .D(
        \mem[27][1] ), .S0(n822), .S1(n828), .Y(n687) );
  MXI4X1 U588 ( .A(n639), .B(n637), .C(n638), .D(n636), .S0(n850), .S1(n843), 
        .Y(n780) );
  MX4X1 U589 ( .A(\mem[92][2] ), .B(\mem[93][2] ), .C(\mem[94][2] ), .D(
        \mem[95][2] ), .S0(n818), .S1(n838), .Y(n636) );
  MX4X1 U590 ( .A(\mem[84][2] ), .B(\mem[85][2] ), .C(\mem[86][2] ), .D(
        \mem[87][2] ), .S0(n818), .S1(n838), .Y(n638) );
  MX4X1 U591 ( .A(\mem[88][2] ), .B(\mem[89][2] ), .C(\mem[90][2] ), .D(
        \mem[91][2] ), .S0(n818), .S1(n838), .Y(n637) );
  MXI4X1 U592 ( .A(n655), .B(n653), .C(n654), .D(n652), .S0(n850), .S1(n846), 
        .Y(n784) );
  MX4X1 U593 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .C(\mem[30][2] ), .D(
        \mem[31][2] ), .S0(n819), .S1(n839), .Y(n652) );
  MX4X1 U594 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .C(\mem[22][2] ), .D(
        \mem[23][2] ), .S0(n819), .S1(n839), .Y(n654) );
  MX4X1 U595 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .C(\mem[26][2] ), .D(
        \mem[27][2] ), .S0(n819), .S1(n839), .Y(n653) );
  MXI4X1 U596 ( .A(n605), .B(n603), .C(n604), .D(n602), .S0(n849), .S1(n845), 
        .Y(n772) );
  MX4X1 U597 ( .A(\mem[92][3] ), .B(\mem[93][3] ), .C(\mem[94][3] ), .D(
        \mem[95][3] ), .S0(n815), .S1(n835), .Y(n602) );
  MX4X1 U598 ( .A(\mem[84][3] ), .B(\mem[85][3] ), .C(\mem[86][3] ), .D(
        \mem[87][3] ), .S0(n815), .S1(n835), .Y(n604) );
  MX4X1 U599 ( .A(\mem[88][3] ), .B(\mem[89][3] ), .C(\mem[90][3] ), .D(
        \mem[91][3] ), .S0(n815), .S1(n835), .Y(n603) );
  MXI4X1 U600 ( .A(n621), .B(n619), .C(n620), .D(n618), .S0(n849), .S1(n845), 
        .Y(n776) );
  MX4X1 U601 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .C(\mem[30][3] ), .D(
        \mem[31][3] ), .S0(n817), .S1(n837), .Y(n618) );
  MX4X1 U602 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .C(\mem[22][3] ), .D(
        \mem[23][3] ), .S0(n817), .S1(n837), .Y(n620) );
  MX4X1 U603 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .C(\mem[26][3] ), .D(
        \mem[27][3] ), .S0(n817), .S1(n837), .Y(n619) );
  MXI4X1 U604 ( .A(n435), .B(n150), .C(n151), .D(n149), .S0(n850), .S1(n844), 
        .Y(n764) );
  MX4X1 U605 ( .A(\mem[92][4] ), .B(\mem[93][4] ), .C(\mem[94][4] ), .D(
        \mem[95][4] ), .S0(n802), .S1(n828), .Y(n149) );
  MX4X1 U606 ( .A(\mem[84][4] ), .B(\mem[85][4] ), .C(\mem[86][4] ), .D(
        \mem[87][4] ), .S0(n802), .S1(n829), .Y(n151) );
  MX4X1 U607 ( .A(\mem[88][4] ), .B(\mem[89][4] ), .C(\mem[90][4] ), .D(
        \mem[91][4] ), .S0(n804), .S1(n829), .Y(n150) );
  MXI4X1 U608 ( .A(n587), .B(n585), .C(n586), .D(n584), .S0(n849), .S1(n845), 
        .Y(n768) );
  MX4X1 U609 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .C(\mem[30][4] ), .D(
        \mem[31][4] ), .S0(n803), .S1(n834), .Y(n584) );
  MX4X1 U610 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .C(\mem[22][4] ), .D(
        \mem[23][4] ), .S0(n802), .S1(n834), .Y(n586) );
  MX4X1 U611 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .C(\mem[26][4] ), .D(
        \mem[27][4] ), .S0(n804), .S1(n834), .Y(n585) );
  MXI4X1 U612 ( .A(n118), .B(n116), .C(n117), .D(n115), .S0(n847), .S1(n844), 
        .Y(n756) );
  MX4X1 U613 ( .A(\mem[92][5] ), .B(\mem[93][5] ), .C(\mem[94][5] ), .D(
        \mem[95][5] ), .S0(n813), .S1(n837), .Y(n115) );
  MX4X1 U614 ( .A(\mem[84][5] ), .B(\mem[85][5] ), .C(\mem[86][5] ), .D(
        \mem[87][5] ), .S0(n814), .S1(n831), .Y(n117) );
  MX4X1 U615 ( .A(\mem[88][5] ), .B(\mem[89][5] ), .C(\mem[90][5] ), .D(
        \mem[91][5] ), .S0(n813), .S1(n828), .Y(n116) );
  MXI4X1 U616 ( .A(n134), .B(n132), .C(n133), .D(n131), .S0(n847), .S1(n844), 
        .Y(n760) );
  MX4X1 U617 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .C(\mem[30][5] ), .D(
        \mem[31][5] ), .S0(n802), .S1(n828), .Y(n131) );
  MX4X1 U618 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .C(\mem[22][5] ), .D(
        \mem[23][5] ), .S0(n804), .S1(n833), .Y(n133) );
  MX4X1 U619 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .C(\mem[26][5] ), .D(
        \mem[27][5] ), .S0(n803), .S1(n829), .Y(n132) );
  MXI4X1 U620 ( .A(n84), .B(n82), .C(n83), .D(n81), .S0(n849), .S1(n843), .Y(
        n748) );
  MX4X1 U621 ( .A(\mem[92][6] ), .B(\mem[93][6] ), .C(\mem[94][6] ), .D(
        \mem[95][6] ), .S0(n811), .S1(n838), .Y(n81) );
  MX4X1 U622 ( .A(\mem[84][6] ), .B(\mem[85][6] ), .C(\mem[86][6] ), .D(
        \mem[87][6] ), .S0(n811), .S1(n825), .Y(n83) );
  MX4X1 U623 ( .A(\mem[88][6] ), .B(\mem[89][6] ), .C(\mem[90][6] ), .D(
        \mem[91][6] ), .S0(n811), .S1(n833), .Y(n82) );
  MXI4X1 U624 ( .A(n100), .B(n98), .C(n99), .D(n97), .S0(n850), .S1(n843), .Y(
        n752) );
  MX4X1 U625 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .C(\mem[30][6] ), .D(
        \mem[31][6] ), .S0(n812), .S1(n833), .Y(n97) );
  MX4X1 U626 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .C(\mem[22][6] ), .D(
        \mem[23][6] ), .S0(n812), .S1(n833), .Y(n99) );
  MX4X1 U627 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .C(\mem[26][6] ), .D(
        \mem[27][6] ), .S0(n812), .S1(n833), .Y(n98) );
  MXI4X1 U628 ( .A(n50), .B(n48), .C(n49), .D(n47), .S0(n848), .S1(n843), .Y(
        n740) );
  MX4X1 U629 ( .A(\mem[92][7] ), .B(\mem[93][7] ), .C(\mem[94][7] ), .D(
        \mem[95][7] ), .S0(n808), .S1(n841), .Y(n47) );
  MX4X1 U630 ( .A(\mem[84][7] ), .B(\mem[85][7] ), .C(\mem[86][7] ), .D(
        \mem[87][7] ), .S0(n809), .S1(n831), .Y(n49) );
  MX4X1 U631 ( .A(\mem[88][7] ), .B(\mem[89][7] ), .C(\mem[90][7] ), .D(
        \mem[91][7] ), .S0(n809), .S1(n831), .Y(n48) );
  MXI4X1 U632 ( .A(n66), .B(n64), .C(n65), .D(n63), .S0(n847), .S1(n843), .Y(
        n744) );
  MX4X1 U633 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .C(\mem[30][7] ), .D(
        \mem[31][7] ), .S0(n810), .S1(n832), .Y(n63) );
  MX4X1 U634 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .C(\mem[22][7] ), .D(
        \mem[23][7] ), .S0(n810), .S1(n832), .Y(n65) );
  MX4X1 U635 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .C(\mem[26][7] ), .D(
        \mem[27][7] ), .S0(n810), .S1(n832), .Y(n64) );
  MXI4X1 U636 ( .A(n16), .B(n14), .C(n15), .D(n13), .S0(n848), .S1(n846), .Y(
        n732) );
  MX4X1 U637 ( .A(valid_mem[92]), .B(valid_mem[93]), .C(valid_mem[94]), .D(
        valid_mem[95]), .S0(n806), .S1(n830), .Y(n13) );
  MX4X1 U638 ( .A(valid_mem[84]), .B(valid_mem[85]), .C(valid_mem[86]), .D(
        valid_mem[87]), .S0(n806), .S1(n825), .Y(n15) );
  MX4X1 U639 ( .A(valid_mem[88]), .B(valid_mem[89]), .C(valid_mem[90]), .D(
        valid_mem[91]), .S0(n806), .S1(n831), .Y(n14) );
  MXI4X1 U640 ( .A(n32), .B(n30), .C(n31), .D(n29), .S0(n848), .S1(n843), .Y(
        n736) );
  MX4X1 U641 ( .A(valid_mem[28]), .B(valid_mem[29]), .C(valid_mem[30]), .D(
        valid_mem[31]), .S0(n807), .S1(n830), .Y(n29) );
  MX4X1 U642 ( .A(valid_mem[20]), .B(valid_mem[21]), .C(valid_mem[22]), .D(
        valid_mem[23]), .S0(n807), .S1(n830), .Y(n31) );
  MX4X1 U643 ( .A(valid_mem[24]), .B(valid_mem[25]), .C(valid_mem[26]), .D(
        valid_mem[27]), .S0(n807), .S1(n830), .Y(n30) );
  MXI4X1 U644 ( .A(n711), .B(n709), .C(n710), .D(n708), .S0(n851), .S1(n846), 
        .Y(n797) );
  MX4X1 U645 ( .A(\mem[76][0] ), .B(\mem[77][0] ), .C(\mem[78][0] ), .D(
        \mem[79][0] ), .S0(n823), .S1(n827), .Y(n708) );
  MX4X1 U646 ( .A(\mem[68][0] ), .B(\mem[69][0] ), .C(\mem[70][0] ), .D(
        \mem[71][0] ), .S0(n823), .S1(n834), .Y(n710) );
  MX4X1 U647 ( .A(\mem[72][0] ), .B(\mem[73][0] ), .C(\mem[74][0] ), .D(
        \mem[75][0] ), .S0(n823), .S1(n829), .Y(n709) );
  MXI4X1 U648 ( .A(n677), .B(n675), .C(n676), .D(n674), .S0(n850), .S1(n846), 
        .Y(n789) );
  MX4X1 U649 ( .A(\mem[76][1] ), .B(\mem[77][1] ), .C(\mem[78][1] ), .D(
        \mem[79][1] ), .S0(n821), .S1(n841), .Y(n674) );
  MX4X1 U650 ( .A(\mem[68][1] ), .B(\mem[69][1] ), .C(\mem[70][1] ), .D(
        \mem[71][1] ), .S0(n821), .S1(n841), .Y(n676) );
  MX4X1 U651 ( .A(\mem[72][1] ), .B(\mem[73][1] ), .C(\mem[74][1] ), .D(
        \mem[75][1] ), .S0(n821), .S1(n841), .Y(n675) );
  MXI4X1 U652 ( .A(n643), .B(n641), .C(n642), .D(n640), .S0(n850), .S1(n845), 
        .Y(n781) );
  MX4X1 U653 ( .A(\mem[76][2] ), .B(\mem[77][2] ), .C(\mem[78][2] ), .D(
        \mem[79][2] ), .S0(n818), .S1(n838), .Y(n640) );
  MX4X1 U654 ( .A(\mem[68][2] ), .B(\mem[69][2] ), .C(\mem[70][2] ), .D(
        \mem[71][2] ), .S0(n818), .S1(n838), .Y(n642) );
  MX4X1 U655 ( .A(\mem[72][2] ), .B(\mem[73][2] ), .C(\mem[74][2] ), .D(
        \mem[75][2] ), .S0(n818), .S1(n838), .Y(n641) );
  MXI4X1 U656 ( .A(n609), .B(n607), .C(n608), .D(n606), .S0(n849), .S1(n845), 
        .Y(n773) );
  MX4X1 U657 ( .A(\mem[76][3] ), .B(\mem[77][3] ), .C(\mem[78][3] ), .D(
        \mem[79][3] ), .S0(n816), .S1(n836), .Y(n606) );
  MX4X1 U658 ( .A(\mem[68][3] ), .B(\mem[69][3] ), .C(\mem[70][3] ), .D(
        \mem[71][3] ), .S0(n816), .S1(n836), .Y(n608) );
  MX4X1 U659 ( .A(\mem[72][3] ), .B(\mem[73][3] ), .C(\mem[74][3] ), .D(
        \mem[75][3] ), .S0(n816), .S1(n836), .Y(n607) );
  MXI4X1 U660 ( .A(n439), .B(n437), .C(n438), .D(n436), .S0(n847), .S1(n844), 
        .Y(n765) );
  MX4X1 U661 ( .A(\mem[76][4] ), .B(\mem[77][4] ), .C(\mem[78][4] ), .D(
        \mem[79][4] ), .S0(n805), .S1(n825), .Y(n436) );
  MX4X1 U662 ( .A(\mem[68][4] ), .B(\mem[69][4] ), .C(\mem[70][4] ), .D(
        \mem[71][4] ), .S0(n805), .S1(n826), .Y(n438) );
  MX4X1 U663 ( .A(\mem[72][4] ), .B(\mem[73][4] ), .C(\mem[74][4] ), .D(
        \mem[75][4] ), .S0(n805), .S1(n826), .Y(n437) );
  MXI4X1 U664 ( .A(n122), .B(n120), .C(n121), .D(n119), .S0(n848), .S1(n844), 
        .Y(n757) );
  MX4X1 U665 ( .A(\mem[76][5] ), .B(\mem[77][5] ), .C(\mem[78][5] ), .D(
        \mem[79][5] ), .S0(n814), .S1(n828), .Y(n119) );
  MX4X1 U666 ( .A(\mem[68][5] ), .B(\mem[69][5] ), .C(\mem[70][5] ), .D(
        \mem[71][5] ), .S0(n814), .S1(n827), .Y(n121) );
  MX4X1 U667 ( .A(\mem[72][5] ), .B(\mem[73][5] ), .C(\mem[74][5] ), .D(
        \mem[75][5] ), .S0(n814), .S1(n841), .Y(n120) );
  MXI4X1 U668 ( .A(n88), .B(n86), .C(n87), .D(n85), .S0(n847), .S1(n843), .Y(
        n749) );
  MX4X1 U669 ( .A(\mem[76][6] ), .B(\mem[77][6] ), .C(\mem[78][6] ), .D(
        \mem[79][6] ), .S0(n811), .S1(n828), .Y(n85) );
  MX4X1 U670 ( .A(\mem[68][6] ), .B(\mem[69][6] ), .C(\mem[70][6] ), .D(
        \mem[71][6] ), .S0(n811), .S1(n826), .Y(n87) );
  MX4X1 U671 ( .A(\mem[72][6] ), .B(\mem[73][6] ), .C(\mem[74][6] ), .D(
        \mem[75][6] ), .S0(n811), .S1(n827), .Y(n86) );
  MXI4X1 U672 ( .A(n54), .B(n52), .C(n53), .D(n51), .S0(n848), .S1(N28), .Y(
        n741) );
  MX4X1 U673 ( .A(\mem[76][7] ), .B(\mem[77][7] ), .C(\mem[78][7] ), .D(
        \mem[79][7] ), .S0(n809), .S1(n831), .Y(n51) );
  MX4X1 U674 ( .A(\mem[68][7] ), .B(\mem[69][7] ), .C(\mem[70][7] ), .D(
        \mem[71][7] ), .S0(n809), .S1(n831), .Y(n53) );
  MX4X1 U675 ( .A(\mem[72][7] ), .B(\mem[73][7] ), .C(\mem[74][7] ), .D(
        \mem[75][7] ), .S0(n809), .S1(n831), .Y(n52) );
  MXI4X1 U676 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n848), .S1(n843), .Y(
        n733) );
  MX4X1 U677 ( .A(valid_mem[76]), .B(valid_mem[77]), .C(valid_mem[78]), .D(
        valid_mem[79]), .S0(n806), .S1(n836), .Y(n17) );
  MX4X1 U678 ( .A(valid_mem[68]), .B(valid_mem[69]), .C(valid_mem[70]), .D(
        valid_mem[71]), .S0(n806), .S1(n827), .Y(n19) );
  MX4X1 U679 ( .A(valid_mem[72]), .B(valid_mem[73]), .C(valid_mem[74]), .D(
        valid_mem[75]), .S0(n806), .S1(n834), .Y(n18) );
  MXI4X1 U680 ( .A(n699), .B(n697), .C(n698), .D(n696), .S0(n851), .S1(n846), 
        .Y(n794) );
  MX4X1 U681 ( .A(\mem[124][0] ), .B(\mem[125][0] ), .C(\mem[126][0] ), .D(
        \mem[127][0] ), .S0(n822), .S1(n827), .Y(n696) );
  MX4X1 U682 ( .A(\mem[116][0] ), .B(\mem[117][0] ), .C(\mem[118][0] ), .D(
        \mem[119][0] ), .S0(n822), .S1(n830), .Y(n698) );
  MX4X1 U683 ( .A(\mem[120][0] ), .B(\mem[121][0] ), .C(\mem[122][0] ), .D(
        \mem[123][0] ), .S0(n822), .S1(n826), .Y(n697) );
  MXI4X1 U684 ( .A(n715), .B(n713), .C(n714), .D(n712), .S0(n851), .S1(n846), 
        .Y(n798) );
  MX4X1 U685 ( .A(\mem[60][0] ), .B(\mem[61][0] ), .C(\mem[62][0] ), .D(
        \mem[63][0] ), .S0(n823), .S1(n829), .Y(n712) );
  MX4X1 U686 ( .A(\mem[52][0] ), .B(\mem[53][0] ), .C(\mem[54][0] ), .D(
        \mem[55][0] ), .S0(n823), .S1(n829), .Y(n714) );
  MX4X1 U687 ( .A(\mem[48][0] ), .B(\mem[49][0] ), .C(\mem[50][0] ), .D(
        \mem[51][0] ), .S0(n824), .S1(n842), .Y(n715) );
  MXI4X1 U688 ( .A(n665), .B(n663), .C(n664), .D(n662), .S0(n850), .S1(n845), 
        .Y(n786) );
  MX4X1 U689 ( .A(\mem[124][1] ), .B(\mem[125][1] ), .C(\mem[126][1] ), .D(
        \mem[127][1] ), .S0(n820), .S1(n840), .Y(n662) );
  MX4X1 U690 ( .A(\mem[116][1] ), .B(\mem[117][1] ), .C(\mem[118][1] ), .D(
        \mem[119][1] ), .S0(n820), .S1(n840), .Y(n664) );
  MX4X1 U691 ( .A(\mem[120][1] ), .B(\mem[121][1] ), .C(\mem[122][1] ), .D(
        \mem[123][1] ), .S0(n820), .S1(n840), .Y(n663) );
  MXI4X1 U692 ( .A(n681), .B(n679), .C(n680), .D(n678), .S0(n851), .S1(n846), 
        .Y(n790) );
  MX4X1 U693 ( .A(\mem[60][1] ), .B(\mem[61][1] ), .C(\mem[62][1] ), .D(
        \mem[63][1] ), .S0(n821), .S1(n841), .Y(n678) );
  MX4X1 U694 ( .A(\mem[52][1] ), .B(\mem[53][1] ), .C(\mem[54][1] ), .D(
        \mem[55][1] ), .S0(n821), .S1(n841), .Y(n680) );
  MX4X1 U695 ( .A(\mem[56][1] ), .B(\mem[57][1] ), .C(\mem[58][1] ), .D(
        \mem[59][1] ), .S0(n821), .S1(n841), .Y(n679) );
  MXI4X1 U696 ( .A(n631), .B(n629), .C(n630), .D(n628), .S0(n850), .S1(n844), 
        .Y(n778) );
  MX4X1 U697 ( .A(\mem[124][2] ), .B(\mem[125][2] ), .C(\mem[126][2] ), .D(
        \mem[127][2] ), .S0(n817), .S1(n837), .Y(n628) );
  MX4X1 U698 ( .A(\mem[116][2] ), .B(\mem[117][2] ), .C(\mem[118][2] ), .D(
        \mem[119][2] ), .S0(n817), .S1(n837), .Y(n630) );
  MX4X1 U699 ( .A(\mem[120][2] ), .B(\mem[121][2] ), .C(\mem[122][2] ), .D(
        \mem[123][2] ), .S0(n817), .S1(n837), .Y(n629) );
  MXI4X1 U700 ( .A(n647), .B(n645), .C(n646), .D(n644), .S0(n850), .S1(n844), 
        .Y(n782) );
  MX4X1 U701 ( .A(\mem[60][2] ), .B(\mem[61][2] ), .C(\mem[62][2] ), .D(
        \mem[63][2] ), .S0(n818), .S1(n838), .Y(n644) );
  MX4X1 U702 ( .A(\mem[52][2] ), .B(\mem[53][2] ), .C(\mem[54][2] ), .D(
        \mem[55][2] ), .S0(n819), .S1(n839), .Y(n646) );
  MX4X1 U703 ( .A(\mem[56][2] ), .B(\mem[57][2] ), .C(\mem[58][2] ), .D(
        \mem[59][2] ), .S0(n818), .S1(n838), .Y(n645) );
  MXI4X1 U704 ( .A(n597), .B(n595), .C(n596), .D(n594), .S0(n849), .S1(n845), 
        .Y(n770) );
  MX4X1 U705 ( .A(\mem[124][3] ), .B(\mem[125][3] ), .C(\mem[126][3] ), .D(
        \mem[127][3] ), .S0(n815), .S1(n835), .Y(n594) );
  MX4X1 U706 ( .A(\mem[116][3] ), .B(\mem[117][3] ), .C(\mem[118][3] ), .D(
        \mem[119][3] ), .S0(n815), .S1(n835), .Y(n596) );
  MX4X1 U707 ( .A(\mem[120][3] ), .B(\mem[121][3] ), .C(\mem[122][3] ), .D(
        \mem[123][3] ), .S0(n815), .S1(n835), .Y(n595) );
  MXI4X1 U708 ( .A(n613), .B(n611), .C(n612), .D(n610), .S0(n849), .S1(n845), 
        .Y(n774) );
  MX4X1 U709 ( .A(\mem[60][3] ), .B(\mem[61][3] ), .C(\mem[62][3] ), .D(
        \mem[63][3] ), .S0(n816), .S1(n836), .Y(n610) );
  MX4X1 U710 ( .A(\mem[52][3] ), .B(\mem[53][3] ), .C(\mem[54][3] ), .D(
        \mem[55][3] ), .S0(n816), .S1(n836), .Y(n612) );
  MX4X1 U711 ( .A(\mem[56][3] ), .B(\mem[57][3] ), .C(\mem[58][3] ), .D(
        \mem[59][3] ), .S0(n816), .S1(n836), .Y(n611) );
  MXI4X1 U712 ( .A(n144), .B(n142), .C(n143), .D(n141), .S0(n849), .S1(n844), 
        .Y(n762) );
  MX4X1 U713 ( .A(\mem[124][4] ), .B(\mem[125][4] ), .C(\mem[126][4] ), .D(
        \mem[127][4] ), .S0(n803), .S1(n828), .Y(n141) );
  MX4X1 U714 ( .A(\mem[116][4] ), .B(\mem[117][4] ), .C(\mem[118][4] ), .D(
        \mem[119][4] ), .S0(n802), .S1(n825), .Y(n143) );
  MX4X1 U715 ( .A(\mem[120][4] ), .B(\mem[121][4] ), .C(\mem[122][4] ), .D(
        \mem[123][4] ), .S0(n804), .S1(n829), .Y(n142) );
  MXI4X1 U716 ( .A(n579), .B(n577), .C(n578), .D(n576), .S0(n849), .S1(n845), 
        .Y(n766) );
  MX4X1 U717 ( .A(\mem[60][4] ), .B(\mem[61][4] ), .C(\mem[62][4] ), .D(
        \mem[63][4] ), .S0(n802), .S1(n825), .Y(n576) );
  MX4X1 U718 ( .A(\mem[52][4] ), .B(\mem[53][4] ), .C(\mem[54][4] ), .D(
        \mem[55][4] ), .S0(n804), .S1(n834), .Y(n578) );
  MX4X1 U719 ( .A(\mem[56][4] ), .B(\mem[57][4] ), .C(\mem[58][4] ), .D(
        \mem[59][4] ), .S0(n803), .S1(n834), .Y(n577) );
  MXI4X1 U720 ( .A(n110), .B(n108), .C(n109), .D(n107), .S0(n851), .S1(n844), 
        .Y(n754) );
  MX4X1 U721 ( .A(\mem[124][5] ), .B(\mem[125][5] ), .C(\mem[126][5] ), .D(
        \mem[127][5] ), .S0(n813), .S1(n829), .Y(n107) );
  MX4X1 U722 ( .A(\mem[116][5] ), .B(\mem[117][5] ), .C(\mem[118][5] ), .D(
        \mem[119][5] ), .S0(n813), .S1(n829), .Y(n109) );
  MX4X1 U723 ( .A(\mem[120][5] ), .B(\mem[121][5] ), .C(\mem[122][5] ), .D(
        \mem[123][5] ), .S0(n813), .S1(n839), .Y(n108) );
  MXI4X1 U724 ( .A(n126), .B(n124), .C(n125), .D(n123), .S0(n847), .S1(n844), 
        .Y(n758) );
  MX4X1 U725 ( .A(\mem[60][5] ), .B(\mem[61][5] ), .C(\mem[62][5] ), .D(
        \mem[63][5] ), .S0(n814), .S1(n838), .Y(n123) );
  MX4X1 U726 ( .A(\mem[52][5] ), .B(\mem[53][5] ), .C(\mem[54][5] ), .D(
        \mem[55][5] ), .S0(n814), .S1(n834), .Y(n125) );
  MX4X1 U727 ( .A(\mem[56][5] ), .B(\mem[57][5] ), .C(\mem[58][5] ), .D(
        \mem[59][5] ), .S0(n814), .S1(n837), .Y(n124) );
  MXI4X1 U728 ( .A(n76), .B(n74), .C(n75), .D(n73), .S0(n848), .S1(n843), .Y(
        n746) );
  MX4X1 U729 ( .A(\mem[124][6] ), .B(\mem[125][6] ), .C(\mem[126][6] ), .D(
        \mem[127][6] ), .S0(n810), .S1(n832), .Y(n73) );
  MX4X1 U730 ( .A(\mem[116][6] ), .B(\mem[117][6] ), .C(\mem[118][6] ), .D(
        \mem[119][6] ), .S0(n810), .S1(n832), .Y(n75) );
  MX4X1 U731 ( .A(\mem[120][6] ), .B(\mem[121][6] ), .C(\mem[122][6] ), .D(
        \mem[123][6] ), .S0(n810), .S1(n832), .Y(n74) );
  MXI4X1 U732 ( .A(n92), .B(n90), .C(n91), .D(n89), .S0(n847), .S1(n843), .Y(
        n750) );
  MX4X1 U733 ( .A(\mem[60][6] ), .B(\mem[61][6] ), .C(\mem[62][6] ), .D(
        \mem[63][6] ), .S0(n812), .S1(n833), .Y(n89) );
  MX4X1 U734 ( .A(\mem[52][6] ), .B(\mem[53][6] ), .C(\mem[54][6] ), .D(
        \mem[55][6] ), .S0(n812), .S1(n833), .Y(n91) );
  MX4X1 U735 ( .A(\mem[56][6] ), .B(\mem[57][6] ), .C(\mem[58][6] ), .D(
        \mem[59][6] ), .S0(n812), .S1(n833), .Y(n90) );
  MXI4X1 U736 ( .A(n42), .B(n40), .C(n41), .D(n39), .S0(n848), .S1(n845), .Y(
        n738) );
  MX4X1 U737 ( .A(\mem[124][7] ), .B(\mem[125][7] ), .C(\mem[126][7] ), .D(
        \mem[127][7] ), .S0(n808), .S1(n841), .Y(n39) );
  MX4X1 U738 ( .A(\mem[116][7] ), .B(\mem[117][7] ), .C(\mem[118][7] ), .D(
        \mem[119][7] ), .S0(n808), .S1(n828), .Y(n41) );
  MX4X1 U739 ( .A(\mem[120][7] ), .B(\mem[121][7] ), .C(\mem[122][7] ), .D(
        \mem[123][7] ), .S0(n808), .S1(n826), .Y(n40) );
  MXI4X1 U740 ( .A(n58), .B(n56), .C(n57), .D(n55), .S0(n851), .S1(n843), .Y(
        n742) );
  MX4X1 U741 ( .A(\mem[60][7] ), .B(\mem[61][7] ), .C(\mem[62][7] ), .D(
        \mem[63][7] ), .S0(n809), .S1(n831), .Y(n55) );
  MX4X1 U742 ( .A(\mem[52][7] ), .B(\mem[53][7] ), .C(\mem[54][7] ), .D(
        \mem[55][7] ), .S0(n809), .S1(n831), .Y(n57) );
  MX4X1 U743 ( .A(\mem[56][7] ), .B(\mem[57][7] ), .C(\mem[58][7] ), .D(
        \mem[59][7] ), .S0(n809), .S1(n831), .Y(n56) );
  MXI4X1 U744 ( .A(n8), .B(n6), .C(n7), .D(n5), .S0(n848), .S1(n844), .Y(n730)
         );
  MX4X1 U745 ( .A(valid_mem[124]), .B(valid_mem[125]), .C(valid_mem[126]), .D(
        valid_mem[127]), .S0(n802), .S1(n827), .Y(n5) );
  MX4X1 U746 ( .A(valid_mem[120]), .B(valid_mem[121]), .C(valid_mem[122]), .D(
        valid_mem[123]), .S0(n805), .S1(n842), .Y(n6) );
  MX4X1 U747 ( .A(valid_mem[116]), .B(valid_mem[117]), .C(valid_mem[118]), .D(
        valid_mem[119]), .S0(n806), .S1(n832), .Y(n7) );
  MXI4X1 U748 ( .A(n24), .B(n22), .C(n23), .D(n21), .S0(n848), .S1(n845), .Y(
        n734) );
  MX4X1 U749 ( .A(valid_mem[60]), .B(valid_mem[61]), .C(valid_mem[62]), .D(
        valid_mem[63]), .S0(n807), .S1(n830), .Y(n21) );
  MX4X1 U750 ( .A(valid_mem[52]), .B(valid_mem[53]), .C(valid_mem[54]), .D(
        valid_mem[55]), .S0(n807), .S1(n830), .Y(n23) );
  MX4X1 U751 ( .A(valid_mem[56]), .B(valid_mem[57]), .C(valid_mem[58]), .D(
        valid_mem[59]), .S0(n807), .S1(n830), .Y(n22) );
  NAND2X1 U752 ( .A(n1475), .B(n1474), .Y(n1193) );
  OAI21XL U753 ( .A0(n869), .A1(n1473), .B0(valid_mem[123]), .Y(n1474) );
  NAND2X1 U754 ( .A(n1472), .B(n1471), .Y(n1192) );
  OAI21XL U755 ( .A0(n869), .A1(n1470), .B0(valid_mem[122]), .Y(n1471) );
  NAND2X1 U756 ( .A(n1469), .B(n1468), .Y(n1191) );
  OAI21XL U757 ( .A0(n869), .A1(n1467), .B0(valid_mem[121]), .Y(n1468) );
  NAND2X1 U758 ( .A(n1466), .B(n1465), .Y(n1190) );
  OAI21XL U759 ( .A0(n869), .A1(n1464), .B0(valid_mem[120]), .Y(n1465) );
  NAND2X1 U760 ( .A(n1463), .B(n1462), .Y(n1189) );
  OAI21XL U761 ( .A0(n869), .A1(n1461), .B0(valid_mem[119]), .Y(n1462) );
  NAND2X1 U762 ( .A(n1460), .B(n1459), .Y(n1188) );
  OAI21XL U763 ( .A0(n869), .A1(n1458), .B0(valid_mem[118]), .Y(n1459) );
  NAND2X1 U764 ( .A(n1457), .B(n1456), .Y(n1187) );
  OAI21XL U765 ( .A0(n869), .A1(n1455), .B0(valid_mem[117]), .Y(n1456) );
  NAND2X1 U766 ( .A(n1454), .B(n1453), .Y(n1186) );
  OAI21XL U767 ( .A0(n869), .A1(n1452), .B0(valid_mem[116]), .Y(n1453) );
  NAND2X1 U768 ( .A(n1451), .B(n1450), .Y(n1185) );
  OAI21XL U769 ( .A0(n869), .A1(n1449), .B0(valid_mem[115]), .Y(n1450) );
  NAND2X1 U770 ( .A(n1448), .B(n1447), .Y(n1184) );
  OAI21XL U771 ( .A0(n869), .A1(n1446), .B0(valid_mem[114]), .Y(n1447) );
  NAND2X1 U772 ( .A(n1445), .B(n1444), .Y(n1183) );
  OAI21XL U773 ( .A0(n869), .A1(n1443), .B0(valid_mem[113]), .Y(n1444) );
  NAND2X1 U774 ( .A(n1442), .B(n1441), .Y(n1182) );
  OAI21XL U775 ( .A0(n869), .A1(n1440), .B0(valid_mem[112]), .Y(n1441) );
  NAND2X1 U776 ( .A(n1484), .B(n1483), .Y(n1196) );
  OAI21XL U777 ( .A0(n869), .A1(n1482), .B0(valid_mem[126]), .Y(n1483) );
  NAND2X1 U778 ( .A(n1481), .B(n1480), .Y(n1195) );
  OAI21XL U779 ( .A0(n869), .A1(n1479), .B0(valid_mem[125]), .Y(n1480) );
  NAND2X1 U780 ( .A(n1478), .B(n1477), .Y(n1194) );
  OAI21XL U781 ( .A0(n869), .A1(n1476), .B0(valid_mem[124]), .Y(n1477) );
  MXI4X1 U782 ( .A(n703), .B(n701), .C(n702), .D(n700), .S0(n851), .S1(n846), 
        .Y(n795) );
  MX4X1 U783 ( .A(\mem[108][0] ), .B(\mem[109][0] ), .C(\mem[110][0] ), .D(
        \mem[111][0] ), .S0(n822), .S1(n829), .Y(n700) );
  MX4X1 U784 ( .A(\mem[100][0] ), .B(\mem[101][0] ), .C(\mem[102][0] ), .D(
        \mem[103][0] ), .S0(n823), .S1(n828), .Y(n702) );
  MX4X1 U785 ( .A(\mem[104][0] ), .B(\mem[105][0] ), .C(\mem[106][0] ), .D(
        \mem[107][0] ), .S0(n822), .S1(n827), .Y(n701) );
  MXI4X1 U786 ( .A(n719), .B(n717), .C(n718), .D(n716), .S0(n851), .S1(n846), 
        .Y(n799) );
  MX4X1 U787 ( .A(\mem[44][0] ), .B(\mem[45][0] ), .C(\mem[46][0] ), .D(
        \mem[47][0] ), .S0(n824), .S1(n842), .Y(n716) );
  MX4X1 U788 ( .A(\mem[36][0] ), .B(\mem[37][0] ), .C(\mem[38][0] ), .D(
        \mem[39][0] ), .S0(n824), .S1(n842), .Y(n718) );
  MX4X1 U789 ( .A(\mem[40][0] ), .B(\mem[41][0] ), .C(\mem[42][0] ), .D(
        \mem[43][0] ), .S0(n824), .S1(n842), .Y(n717) );
  MXI4X1 U790 ( .A(n669), .B(n667), .C(n668), .D(n666), .S0(n850), .S1(n845), 
        .Y(n787) );
  MX4X1 U791 ( .A(\mem[108][1] ), .B(\mem[109][1] ), .C(\mem[110][1] ), .D(
        \mem[111][1] ), .S0(n820), .S1(n840), .Y(n666) );
  MX4X1 U792 ( .A(\mem[100][1] ), .B(\mem[101][1] ), .C(\mem[102][1] ), .D(
        \mem[103][1] ), .S0(n820), .S1(n840), .Y(n668) );
  MX4X1 U793 ( .A(\mem[104][1] ), .B(\mem[105][1] ), .C(\mem[106][1] ), .D(
        \mem[107][1] ), .S0(n820), .S1(n840), .Y(n667) );
  MXI4X1 U794 ( .A(n685), .B(n683), .C(n684), .D(n682), .S0(n851), .S1(n846), 
        .Y(n791) );
  MX4X1 U795 ( .A(\mem[44][1] ), .B(\mem[45][1] ), .C(\mem[46][1] ), .D(
        \mem[47][1] ), .S0(n821), .S1(n841), .Y(n682) );
  MX4X1 U796 ( .A(\mem[36][1] ), .B(\mem[37][1] ), .C(\mem[38][1] ), .D(
        \mem[39][1] ), .S0(n821), .S1(n841), .Y(n684) );
  MX4X1 U797 ( .A(\mem[40][1] ), .B(\mem[41][1] ), .C(\mem[42][1] ), .D(
        \mem[43][1] ), .S0(n821), .S1(n841), .Y(n683) );
  MXI4X1 U798 ( .A(n635), .B(n633), .C(n634), .D(n632), .S0(n850), .S1(n844), 
        .Y(n779) );
  MX4X1 U799 ( .A(\mem[108][2] ), .B(\mem[109][2] ), .C(\mem[110][2] ), .D(
        \mem[111][2] ), .S0(n817), .S1(n837), .Y(n632) );
  MX4X1 U800 ( .A(\mem[100][2] ), .B(\mem[101][2] ), .C(\mem[102][2] ), .D(
        \mem[103][2] ), .S0(n818), .S1(n838), .Y(n634) );
  MX4X1 U801 ( .A(\mem[104][2] ), .B(\mem[105][2] ), .C(\mem[106][2] ), .D(
        \mem[107][2] ), .S0(n818), .S1(n838), .Y(n633) );
  MXI4X1 U802 ( .A(n651), .B(n649), .C(n650), .D(n648), .S0(n850), .S1(n844), 
        .Y(n783) );
  MX4X1 U803 ( .A(\mem[44][2] ), .B(\mem[45][2] ), .C(\mem[46][2] ), .D(
        \mem[47][2] ), .S0(n819), .S1(n839), .Y(n648) );
  MX4X1 U804 ( .A(\mem[36][2] ), .B(\mem[37][2] ), .C(\mem[38][2] ), .D(
        \mem[39][2] ), .S0(n819), .S1(n839), .Y(n650) );
  MX4X1 U805 ( .A(\mem[40][2] ), .B(\mem[41][2] ), .C(\mem[42][2] ), .D(
        \mem[43][2] ), .S0(n819), .S1(n839), .Y(n649) );
  MXI4X1 U806 ( .A(n601), .B(n599), .C(n600), .D(n598), .S0(n849), .S1(n845), 
        .Y(n771) );
  MX4X1 U807 ( .A(\mem[108][3] ), .B(\mem[109][3] ), .C(\mem[110][3] ), .D(
        \mem[111][3] ), .S0(n815), .S1(n835), .Y(n598) );
  MX4X1 U808 ( .A(\mem[100][3] ), .B(\mem[101][3] ), .C(\mem[102][3] ), .D(
        \mem[103][3] ), .S0(n815), .S1(n835), .Y(n600) );
  MX4X1 U809 ( .A(\mem[104][3] ), .B(\mem[105][3] ), .C(\mem[106][3] ), .D(
        \mem[107][3] ), .S0(n815), .S1(n835), .Y(n599) );
  MXI4X1 U810 ( .A(n617), .B(n615), .C(n616), .D(n614), .S0(n849), .S1(n845), 
        .Y(n775) );
  MX4X1 U811 ( .A(\mem[44][3] ), .B(\mem[45][3] ), .C(\mem[46][3] ), .D(
        \mem[47][3] ), .S0(n816), .S1(n836), .Y(n614) );
  MX4X1 U812 ( .A(\mem[36][3] ), .B(\mem[37][3] ), .C(\mem[38][3] ), .D(
        \mem[39][3] ), .S0(n816), .S1(n836), .Y(n616) );
  MX4X1 U813 ( .A(\mem[40][3] ), .B(\mem[41][3] ), .C(\mem[42][3] ), .D(
        \mem[43][3] ), .S0(n816), .S1(n836), .Y(n615) );
  MXI4X1 U814 ( .A(n148), .B(n146), .C(n147), .D(n145), .S0(n847), .S1(n844), 
        .Y(n763) );
  MX4X1 U815 ( .A(\mem[108][4] ), .B(\mem[109][4] ), .C(\mem[110][4] ), .D(
        \mem[111][4] ), .S0(n805), .S1(n825), .Y(n145) );
  MX4X1 U816 ( .A(\mem[100][4] ), .B(\mem[101][4] ), .C(\mem[102][4] ), .D(
        \mem[103][4] ), .S0(n805), .S1(n826), .Y(n147) );
  MX4X1 U817 ( .A(\mem[104][4] ), .B(\mem[105][4] ), .C(\mem[106][4] ), .D(
        \mem[107][4] ), .S0(n805), .S1(n825), .Y(n146) );
  MXI4X1 U818 ( .A(n583), .B(n581), .C(n582), .D(n580), .S0(n849), .S1(n845), 
        .Y(n767) );
  MX4X1 U819 ( .A(\mem[44][4] ), .B(\mem[45][4] ), .C(\mem[46][4] ), .D(
        \mem[47][4] ), .S0(n802), .S1(n834), .Y(n580) );
  MX4X1 U820 ( .A(\mem[36][4] ), .B(\mem[37][4] ), .C(\mem[38][4] ), .D(
        \mem[39][4] ), .S0(n803), .S1(n834), .Y(n582) );
  MX4X1 U821 ( .A(\mem[40][4] ), .B(\mem[41][4] ), .C(\mem[42][4] ), .D(
        \mem[43][4] ), .S0(n804), .S1(n834), .Y(n581) );
  MXI4X1 U822 ( .A(n114), .B(n112), .C(n113), .D(n111), .S0(n847), .S1(n844), 
        .Y(n755) );
  MX4X1 U823 ( .A(\mem[108][5] ), .B(\mem[109][5] ), .C(\mem[110][5] ), .D(
        \mem[111][5] ), .S0(n813), .S1(n842), .Y(n111) );
  MX4X1 U824 ( .A(\mem[100][5] ), .B(\mem[101][5] ), .C(\mem[102][5] ), .D(
        \mem[103][5] ), .S0(n813), .S1(n834), .Y(n113) );
  MX4X1 U825 ( .A(\mem[104][5] ), .B(\mem[105][5] ), .C(\mem[106][5] ), .D(
        \mem[107][5] ), .S0(n813), .S1(n826), .Y(n112) );
  MXI4X1 U826 ( .A(n130), .B(n128), .C(n129), .D(n127), .S0(n850), .S1(n844), 
        .Y(n759) );
  MX4X1 U827 ( .A(\mem[44][5] ), .B(\mem[45][5] ), .C(\mem[46][5] ), .D(
        \mem[47][5] ), .S0(n814), .S1(n842), .Y(n127) );
  MX4X1 U828 ( .A(\mem[36][5] ), .B(\mem[37][5] ), .C(\mem[38][5] ), .D(
        \mem[39][5] ), .S0(n814), .S1(n825), .Y(n129) );
  MX4X1 U829 ( .A(\mem[40][5] ), .B(\mem[41][5] ), .C(\mem[42][5] ), .D(
        \mem[43][5] ), .S0(n814), .S1(n835), .Y(n128) );
  MXI4X1 U830 ( .A(n80), .B(n78), .C(n79), .D(n77), .S0(n847), .S1(n843), .Y(
        n747) );
  MX4X1 U831 ( .A(\mem[108][6] ), .B(\mem[109][6] ), .C(\mem[110][6] ), .D(
        \mem[111][6] ), .S0(n811), .S1(n828), .Y(n77) );
  MX4X1 U832 ( .A(\mem[100][6] ), .B(\mem[101][6] ), .C(\mem[102][6] ), .D(
        \mem[103][6] ), .S0(n811), .S1(n829), .Y(n79) );
  MX4X1 U833 ( .A(\mem[104][6] ), .B(\mem[105][6] ), .C(\mem[106][6] ), .D(
        \mem[107][6] ), .S0(n811), .S1(n827), .Y(n78) );
  MXI4X1 U834 ( .A(n96), .B(n94), .C(n95), .D(n93), .S0(N29), .S1(n843), .Y(
        n751) );
  MX4X1 U835 ( .A(\mem[44][6] ), .B(\mem[45][6] ), .C(\mem[46][6] ), .D(
        \mem[47][6] ), .S0(n812), .S1(n833), .Y(n93) );
  MX4X1 U836 ( .A(\mem[36][6] ), .B(\mem[37][6] ), .C(\mem[38][6] ), .D(
        \mem[39][6] ), .S0(n812), .S1(n833), .Y(n95) );
  MX4X1 U837 ( .A(\mem[40][6] ), .B(\mem[41][6] ), .C(\mem[42][6] ), .D(
        \mem[43][6] ), .S0(n812), .S1(n833), .Y(n94) );
  MXI4X1 U838 ( .A(n46), .B(n44), .C(n45), .D(n43), .S0(n848), .S1(n843), .Y(
        n739) );
  MX4X1 U839 ( .A(\mem[108][7] ), .B(\mem[109][7] ), .C(\mem[110][7] ), .D(
        \mem[111][7] ), .S0(n808), .S1(n831), .Y(n43) );
  MX4X1 U840 ( .A(\mem[100][7] ), .B(\mem[101][7] ), .C(\mem[102][7] ), .D(
        \mem[103][7] ), .S0(n808), .S1(n839), .Y(n45) );
  MX4X1 U841 ( .A(\mem[104][7] ), .B(\mem[105][7] ), .C(\mem[106][7] ), .D(
        \mem[107][7] ), .S0(n808), .S1(n835), .Y(n44) );
  MXI4X1 U842 ( .A(n62), .B(n60), .C(n61), .D(n59), .S0(n847), .S1(n845), .Y(
        n743) );
  MX4X1 U843 ( .A(\mem[44][7] ), .B(\mem[45][7] ), .C(\mem[46][7] ), .D(
        \mem[47][7] ), .S0(n809), .S1(n831), .Y(n59) );
  MX4X1 U844 ( .A(\mem[36][7] ), .B(\mem[37][7] ), .C(\mem[38][7] ), .D(
        \mem[39][7] ), .S0(n810), .S1(n832), .Y(n61) );
  MX4X1 U845 ( .A(\mem[40][7] ), .B(\mem[41][7] ), .C(\mem[42][7] ), .D(
        \mem[43][7] ), .S0(n809), .S1(n831), .Y(n60) );
  MXI4X1 U846 ( .A(n12), .B(n10), .C(n11), .D(n9), .S0(n848), .S1(n843), .Y(
        n731) );
  MX4X1 U847 ( .A(valid_mem[108]), .B(valid_mem[109]), .C(valid_mem[110]), .D(
        valid_mem[111]), .S0(n806), .S1(n836), .Y(n9) );
  MX4X1 U848 ( .A(valid_mem[100]), .B(valid_mem[101]), .C(valid_mem[102]), .D(
        valid_mem[103]), .S0(n806), .S1(n833), .Y(n11) );
  MX4X1 U849 ( .A(valid_mem[104]), .B(valid_mem[105]), .C(valid_mem[106]), .D(
        valid_mem[107]), .S0(n806), .S1(n841), .Y(n10) );
  MXI4X1 U850 ( .A(n28), .B(n26), .C(n27), .D(n25), .S0(n848), .S1(n843), .Y(
        n735) );
  MX4X1 U851 ( .A(valid_mem[44]), .B(valid_mem[45]), .C(valid_mem[46]), .D(
        valid_mem[47]), .S0(n807), .S1(n830), .Y(n25) );
  MX4X1 U852 ( .A(valid_mem[36]), .B(valid_mem[37]), .C(valid_mem[38]), .D(
        valid_mem[39]), .S0(n807), .S1(n830), .Y(n27) );
  MX4X1 U853 ( .A(valid_mem[40]), .B(valid_mem[41]), .C(valid_mem[42]), .D(
        valid_mem[43]), .S0(n807), .S1(n830), .Y(n26) );
  NAND2X1 U854 ( .A(n1488), .B(n1487), .Y(n1197) );
  OAI21XL U855 ( .A0(n869), .A1(n1485), .B0(valid_mem[127]), .Y(n1487) );
  NAND2X1 U856 ( .A(n1428), .B(n1427), .Y(n1176) );
  OAI21XL U857 ( .A0(n1470), .A1(n867), .B0(valid_mem[106]), .Y(n1427) );
  NAND2X1 U858 ( .A(n1420), .B(n1419), .Y(n1172) );
  OAI21XL U859 ( .A0(n1458), .A1(n867), .B0(valid_mem[102]), .Y(n1419) );
  NAND2X1 U860 ( .A(n1418), .B(n1417), .Y(n1171) );
  OAI21XL U861 ( .A0(n1455), .A1(n867), .B0(valid_mem[101]), .Y(n1417) );
  NAND2X1 U862 ( .A(n1416), .B(n1415), .Y(n1170) );
  OAI21XL U863 ( .A0(n1452), .A1(n867), .B0(valid_mem[100]), .Y(n1415) );
  NAND2X1 U864 ( .A(n1412), .B(n1411), .Y(n1168) );
  OAI21XL U865 ( .A0(n1446), .A1(n867), .B0(valid_mem[98]), .Y(n1411) );
  NAND2X1 U866 ( .A(n1395), .B(n1394), .Y(n1160) );
  OAI21XL U867 ( .A0(n1470), .A1(n865), .B0(valid_mem[90]), .Y(n1394) );
  NAND2X1 U868 ( .A(n1387), .B(n1386), .Y(n1156) );
  OAI21XL U869 ( .A0(n1458), .A1(n865), .B0(valid_mem[86]), .Y(n1386) );
  NAND2X1 U870 ( .A(n1354), .B(n1353), .Y(n1140) );
  OAI21XL U871 ( .A0(n1458), .A1(n863), .B0(valid_mem[70]), .Y(n1353) );
  NAND2X1 U872 ( .A(n1296), .B(n1295), .Y(n1112) );
  OAI21XL U873 ( .A0(n1470), .A1(n859), .B0(valid_mem[42]), .Y(n1295) );
  NAND2X1 U874 ( .A(n1439), .B(n1438), .Y(n1181) );
  OAI21XL U875 ( .A0(n1485), .A1(n867), .B0(valid_mem[111]), .Y(n1438) );
  NAND2X1 U876 ( .A(n1436), .B(n1435), .Y(n1180) );
  OAI21XL U877 ( .A0(n1482), .A1(n867), .B0(valid_mem[110]), .Y(n1435) );
  NAND2X1 U878 ( .A(n1434), .B(n1433), .Y(n1179) );
  OAI21XL U879 ( .A0(n1479), .A1(n867), .B0(valid_mem[109]), .Y(n1433) );
  NAND2X1 U880 ( .A(n1432), .B(n1431), .Y(n1178) );
  OAI21XL U881 ( .A0(n1476), .A1(n867), .B0(valid_mem[108]), .Y(n1431) );
  NAND2X1 U882 ( .A(n1430), .B(n1429), .Y(n1177) );
  OAI21XL U883 ( .A0(n1473), .A1(n867), .B0(valid_mem[107]), .Y(n1429) );
  NAND2X1 U884 ( .A(n1426), .B(n1425), .Y(n1175) );
  OAI21XL U885 ( .A0(n1467), .A1(n867), .B0(valid_mem[105]), .Y(n1425) );
  NAND2X1 U886 ( .A(n1424), .B(n1423), .Y(n1174) );
  OAI21XL U887 ( .A0(n1464), .A1(n867), .B0(valid_mem[104]), .Y(n1423) );
  NAND2X1 U888 ( .A(n1422), .B(n1421), .Y(n1173) );
  OAI21XL U889 ( .A0(n1461), .A1(n867), .B0(valid_mem[103]), .Y(n1421) );
  NAND2X1 U890 ( .A(n1414), .B(n1413), .Y(n1169) );
  OAI21XL U891 ( .A0(n1449), .A1(n867), .B0(valid_mem[99]), .Y(n1413) );
  NAND2X1 U892 ( .A(n1410), .B(n1409), .Y(n1167) );
  OAI21XL U893 ( .A0(n1443), .A1(n867), .B0(valid_mem[97]), .Y(n1409) );
  NAND2X1 U894 ( .A(n1408), .B(n1407), .Y(n1166) );
  OAI21XL U895 ( .A0(n1440), .A1(n867), .B0(valid_mem[96]), .Y(n1407) );
  NAND2X1 U896 ( .A(n1401), .B(n1400), .Y(n1163) );
  OAI21XL U897 ( .A0(n1479), .A1(n865), .B0(valid_mem[93]), .Y(n1400) );
  NAND2X1 U898 ( .A(n1399), .B(n1398), .Y(n1162) );
  OAI21XL U899 ( .A0(n1476), .A1(n865), .B0(valid_mem[92]), .Y(n1398) );
  NAND2X1 U900 ( .A(n1397), .B(n1396), .Y(n1161) );
  OAI21XL U901 ( .A0(n1473), .A1(n865), .B0(valid_mem[91]), .Y(n1396) );
  NAND2X1 U902 ( .A(n1393), .B(n1392), .Y(n1159) );
  OAI21XL U903 ( .A0(n1467), .A1(n865), .B0(valid_mem[89]), .Y(n1392) );
  NAND2X1 U904 ( .A(n1391), .B(n1390), .Y(n1158) );
  OAI21XL U905 ( .A0(n1464), .A1(n865), .B0(valid_mem[88]), .Y(n1390) );
  NAND2X1 U906 ( .A(n1385), .B(n1384), .Y(n1155) );
  OAI21XL U907 ( .A0(n1455), .A1(n865), .B0(valid_mem[85]), .Y(n1384) );
  NAND2X1 U908 ( .A(n1383), .B(n1382), .Y(n1154) );
  OAI21XL U909 ( .A0(n1452), .A1(n865), .B0(valid_mem[84]), .Y(n1382) );
  NAND2X1 U910 ( .A(n1379), .B(n1378), .Y(n1152) );
  OAI21XL U911 ( .A0(n1446), .A1(n865), .B0(valid_mem[82]), .Y(n1378) );
  NAND2X1 U912 ( .A(n1362), .B(n1361), .Y(n1144) );
  OAI21XL U913 ( .A0(n1470), .A1(n863), .B0(valid_mem[74]), .Y(n1361) );
  NAND2X1 U914 ( .A(n1381), .B(n1380), .Y(n1153) );
  OAI21XL U915 ( .A0(n1449), .A1(n865), .B0(valid_mem[83]), .Y(n1380) );
  NAND2X1 U916 ( .A(n1377), .B(n1376), .Y(n1151) );
  OAI21XL U917 ( .A0(n1443), .A1(n865), .B0(valid_mem[81]), .Y(n1376) );
  NAND2X1 U918 ( .A(n1375), .B(n1374), .Y(n1150) );
  OAI21XL U919 ( .A0(n1440), .A1(n865), .B0(valid_mem[80]), .Y(n1374) );
  NAND2X1 U920 ( .A(n1373), .B(n1372), .Y(n1149) );
  OAI21XL U921 ( .A0(n1485), .A1(n863), .B0(valid_mem[79]), .Y(n1372) );
  NAND2X1 U922 ( .A(n1370), .B(n1369), .Y(n1148) );
  OAI21XL U923 ( .A0(n1482), .A1(n863), .B0(valid_mem[78]), .Y(n1369) );
  NAND2X1 U924 ( .A(n1368), .B(n1367), .Y(n1147) );
  OAI21XL U925 ( .A0(n1479), .A1(n863), .B0(valid_mem[77]), .Y(n1367) );
  NAND2X1 U926 ( .A(n1366), .B(n1365), .Y(n1146) );
  OAI21XL U927 ( .A0(n1476), .A1(n863), .B0(valid_mem[76]), .Y(n1365) );
  NAND2X1 U928 ( .A(n1364), .B(n1363), .Y(n1145) );
  OAI21XL U929 ( .A0(n1473), .A1(n863), .B0(valid_mem[75]), .Y(n1363) );
  NAND2X1 U930 ( .A(n1360), .B(n1359), .Y(n1143) );
  OAI21XL U931 ( .A0(n1467), .A1(n863), .B0(valid_mem[73]), .Y(n1359) );
  NAND2X1 U932 ( .A(n1358), .B(n1357), .Y(n1142) );
  OAI21XL U933 ( .A0(n1464), .A1(n863), .B0(valid_mem[72]), .Y(n1357) );
  NAND2X1 U934 ( .A(n1352), .B(n1351), .Y(n1139) );
  OAI21XL U935 ( .A0(n1455), .A1(n863), .B0(valid_mem[69]), .Y(n1351) );
  NAND2X1 U936 ( .A(n1350), .B(n1349), .Y(n1138) );
  OAI21XL U937 ( .A0(n1452), .A1(n863), .B0(valid_mem[68]), .Y(n1349) );
  NAND2X1 U938 ( .A(n1346), .B(n1345), .Y(n1136) );
  OAI21XL U939 ( .A0(n1446), .A1(n863), .B0(valid_mem[66]), .Y(n1345) );
  NAND2X1 U940 ( .A(n1342), .B(n1341), .Y(n1134) );
  OAI21XL U941 ( .A0(n1440), .A1(n863), .B0(valid_mem[64]), .Y(n1341) );
  NAND2X1 U942 ( .A(n1329), .B(n1328), .Y(n1128) );
  OAI21XL U943 ( .A0(n1470), .A1(n861), .B0(valid_mem[58]), .Y(n1328) );
  NAND2X1 U944 ( .A(n1325), .B(n1324), .Y(n1126) );
  OAI21XL U945 ( .A0(n1464), .A1(n861), .B0(valid_mem[56]), .Y(n1324) );
  NAND2X1 U946 ( .A(n1321), .B(n1320), .Y(n1124) );
  OAI21XL U947 ( .A0(n1458), .A1(n861), .B0(valid_mem[54]), .Y(n1320) );
  NAND2X1 U948 ( .A(n1319), .B(n1318), .Y(n1123) );
  OAI21XL U949 ( .A0(n1455), .A1(n861), .B0(valid_mem[53]), .Y(n1318) );
  NAND2X1 U950 ( .A(n1317), .B(n1316), .Y(n1122) );
  OAI21XL U951 ( .A0(n1452), .A1(n861), .B0(valid_mem[52]), .Y(n1316) );
  NAND2X1 U952 ( .A(n1313), .B(n1312), .Y(n1120) );
  OAI21XL U953 ( .A0(n1446), .A1(n861), .B0(valid_mem[50]), .Y(n1312) );
  NAND2X1 U954 ( .A(n1311), .B(n1310), .Y(n1119) );
  OAI21XL U955 ( .A0(n1443), .A1(n861), .B0(valid_mem[49]), .Y(n1310) );
  NAND2X1 U956 ( .A(n1309), .B(n1308), .Y(n1118) );
  OAI21XL U957 ( .A0(n1440), .A1(n861), .B0(valid_mem[48]), .Y(n1308) );
  NAND2X1 U958 ( .A(n1294), .B(n1293), .Y(n1111) );
  OAI21XL U959 ( .A0(n1467), .A1(n859), .B0(valid_mem[41]), .Y(n1293) );
  NAND2X1 U960 ( .A(n1292), .B(n1291), .Y(n1110) );
  OAI21XL U961 ( .A0(n1464), .A1(n859), .B0(valid_mem[40]), .Y(n1291) );
  NAND2X1 U962 ( .A(n1288), .B(n1287), .Y(n1108) );
  OAI21XL U963 ( .A0(n1458), .A1(n859), .B0(valid_mem[38]), .Y(n1287) );
  NAND2X1 U964 ( .A(n1286), .B(n1285), .Y(n1107) );
  OAI21XL U965 ( .A0(n1455), .A1(n859), .B0(valid_mem[37]), .Y(n1285) );
  NAND2X1 U966 ( .A(n1284), .B(n1283), .Y(n1106) );
  OAI21XL U967 ( .A0(n1452), .A1(n859), .B0(valid_mem[36]), .Y(n1283) );
  NAND2X1 U968 ( .A(n1280), .B(n1279), .Y(n1104) );
  OAI21XL U969 ( .A0(n1446), .A1(n859), .B0(valid_mem[34]), .Y(n1279) );
  NAND2X1 U970 ( .A(n1278), .B(n1277), .Y(n1103) );
  OAI21XL U971 ( .A0(n1443), .A1(n859), .B0(valid_mem[33]), .Y(n1277) );
  NAND2X1 U972 ( .A(n1276), .B(n1275), .Y(n1102) );
  OAI21XL U973 ( .A0(n1440), .A1(n859), .B0(valid_mem[32]), .Y(n1275) );
  NAND2X1 U974 ( .A(n1263), .B(n1262), .Y(n1096) );
  OAI21XL U975 ( .A0(n1470), .A1(n857), .B0(valid_mem[26]), .Y(n1262) );
  NAND2X1 U976 ( .A(n1255), .B(n1254), .Y(n1092) );
  OAI21XL U977 ( .A0(n1458), .A1(n857), .B0(valid_mem[22]), .Y(n1254) );
  NAND2X1 U978 ( .A(n1251), .B(n1250), .Y(n1090) );
  OAI21XL U979 ( .A0(n1452), .A1(n857), .B0(valid_mem[20]), .Y(n1250) );
  NAND2X1 U980 ( .A(n1247), .B(n1246), .Y(n1088) );
  OAI21XL U981 ( .A0(n1446), .A1(n857), .B0(valid_mem[18]), .Y(n1246) );
  NAND2X1 U982 ( .A(n1230), .B(n1229), .Y(n1080) );
  OAI21XL U983 ( .A0(n1470), .A1(n855), .B0(valid_mem[10]), .Y(n1229) );
  NAND2X1 U984 ( .A(n1406), .B(n1405), .Y(n1165) );
  OAI21XL U985 ( .A0(n1485), .A1(n865), .B0(valid_mem[95]), .Y(n1405) );
  NAND2X1 U986 ( .A(n1403), .B(n1402), .Y(n1164) );
  OAI21XL U987 ( .A0(n1482), .A1(n865), .B0(valid_mem[94]), .Y(n1402) );
  NAND2X1 U988 ( .A(n1356), .B(n1355), .Y(n1141) );
  OAI21XL U989 ( .A0(n1461), .A1(n863), .B0(valid_mem[71]), .Y(n1355) );
  NAND2X1 U990 ( .A(n1348), .B(n1347), .Y(n1137) );
  OAI21XL U991 ( .A0(n1449), .A1(n863), .B0(valid_mem[67]), .Y(n1347) );
  NAND2X1 U992 ( .A(n1344), .B(n1343), .Y(n1135) );
  OAI21XL U993 ( .A0(n1443), .A1(n863), .B0(valid_mem[65]), .Y(n1343) );
  NAND2X1 U994 ( .A(n1340), .B(n1339), .Y(n1133) );
  OAI21XL U995 ( .A0(n1485), .A1(n861), .B0(valid_mem[63]), .Y(n1339) );
  NAND2X1 U996 ( .A(n1337), .B(n1336), .Y(n1132) );
  OAI21XL U997 ( .A0(n1482), .A1(n861), .B0(valid_mem[62]), .Y(n1336) );
  NAND2X1 U998 ( .A(n1335), .B(n1334), .Y(n1131) );
  OAI21XL U999 ( .A0(n1479), .A1(n861), .B0(valid_mem[61]), .Y(n1334) );
  NAND2X1 U1000 ( .A(n1333), .B(n1332), .Y(n1130) );
  OAI21XL U1001 ( .A0(n1476), .A1(n861), .B0(valid_mem[60]), .Y(n1332) );
  NAND2X1 U1002 ( .A(n1331), .B(n1330), .Y(n1129) );
  OAI21XL U1003 ( .A0(n1473), .A1(n861), .B0(valid_mem[59]), .Y(n1330) );
  NAND2X1 U1004 ( .A(n1327), .B(n1326), .Y(n1127) );
  OAI21XL U1005 ( .A0(n1467), .A1(n861), .B0(valid_mem[57]), .Y(n1326) );
  NAND2X1 U1006 ( .A(n1323), .B(n1322), .Y(n1125) );
  OAI21XL U1007 ( .A0(n1461), .A1(n861), .B0(valid_mem[55]), .Y(n1322) );
  NAND2X1 U1008 ( .A(n1315), .B(n1314), .Y(n1121) );
  OAI21XL U1009 ( .A0(n1449), .A1(n861), .B0(valid_mem[51]), .Y(n1314) );
  NAND2X1 U1010 ( .A(n1307), .B(n1306), .Y(n1117) );
  OAI21XL U1011 ( .A0(n1485), .A1(n859), .B0(valid_mem[47]), .Y(n1306) );
  NAND2X1 U1012 ( .A(n1304), .B(n1303), .Y(n1116) );
  OAI21XL U1013 ( .A0(n1482), .A1(n859), .B0(valid_mem[46]), .Y(n1303) );
  NAND2X1 U1014 ( .A(n1302), .B(n1301), .Y(n1115) );
  OAI21XL U1015 ( .A0(n1479), .A1(n859), .B0(valid_mem[45]), .Y(n1301) );
  NAND2X1 U1016 ( .A(n1300), .B(n1299), .Y(n1114) );
  OAI21XL U1017 ( .A0(n1476), .A1(n859), .B0(valid_mem[44]), .Y(n1299) );
  NAND2X1 U1018 ( .A(n1298), .B(n1297), .Y(n1113) );
  OAI21XL U1019 ( .A0(n1473), .A1(n859), .B0(valid_mem[43]), .Y(n1297) );
  NAND2X1 U1020 ( .A(n1290), .B(n1289), .Y(n1109) );
  OAI21XL U1021 ( .A0(n1461), .A1(n859), .B0(valid_mem[39]), .Y(n1289) );
  NAND2X1 U1022 ( .A(n1282), .B(n1281), .Y(n1105) );
  OAI21XL U1023 ( .A0(n1449), .A1(n859), .B0(valid_mem[35]), .Y(n1281) );
  NAND2X1 U1024 ( .A(n1274), .B(n1273), .Y(n1101) );
  OAI21XL U1025 ( .A0(n1485), .A1(n857), .B0(valid_mem[31]), .Y(n1273) );
  NAND2X1 U1026 ( .A(n1271), .B(n1270), .Y(n1100) );
  OAI21XL U1027 ( .A0(n1482), .A1(n857), .B0(valid_mem[30]), .Y(n1270) );
  NAND2X1 U1028 ( .A(n1269), .B(n1268), .Y(n1099) );
  OAI21XL U1029 ( .A0(n1479), .A1(n857), .B0(valid_mem[29]), .Y(n1268) );
  NAND2X1 U1030 ( .A(n1267), .B(n1266), .Y(n1098) );
  OAI21XL U1031 ( .A0(n1476), .A1(n857), .B0(valid_mem[28]), .Y(n1266) );
  NAND2X1 U1032 ( .A(n1265), .B(n1264), .Y(n1097) );
  OAI21XL U1033 ( .A0(n1473), .A1(n857), .B0(valid_mem[27]), .Y(n1264) );
  NAND2X1 U1034 ( .A(n1261), .B(n1260), .Y(n1095) );
  OAI21XL U1035 ( .A0(n1467), .A1(n857), .B0(valid_mem[25]), .Y(n1260) );
  NAND2X1 U1036 ( .A(n1259), .B(n1258), .Y(n1094) );
  OAI21XL U1037 ( .A0(n1464), .A1(n857), .B0(valid_mem[24]), .Y(n1258) );
  NAND2X1 U1038 ( .A(n1257), .B(n1256), .Y(n1093) );
  OAI21XL U1039 ( .A0(n1461), .A1(n857), .B0(valid_mem[23]), .Y(n1256) );
  NAND2X1 U1040 ( .A(n1253), .B(n1252), .Y(n1091) );
  OAI21XL U1041 ( .A0(n1455), .A1(n857), .B0(valid_mem[21]), .Y(n1252) );
  NAND2X1 U1042 ( .A(n1249), .B(n1248), .Y(n1089) );
  OAI21XL U1043 ( .A0(n1449), .A1(n857), .B0(valid_mem[19]), .Y(n1248) );
  NAND2X1 U1044 ( .A(n1245), .B(n1244), .Y(n1087) );
  OAI21XL U1045 ( .A0(n1443), .A1(n857), .B0(valid_mem[17]), .Y(n1244) );
  NAND2X1 U1046 ( .A(n1243), .B(n1242), .Y(n1086) );
  OAI21XL U1047 ( .A0(n1440), .A1(n857), .B0(valid_mem[16]), .Y(n1242) );
  NAND2X1 U1048 ( .A(n1241), .B(n1240), .Y(n1085) );
  OAI21XL U1049 ( .A0(n1485), .A1(n855), .B0(valid_mem[15]), .Y(n1240) );
  NAND2X1 U1050 ( .A(n1238), .B(n1237), .Y(n1084) );
  OAI21XL U1051 ( .A0(n1482), .A1(n855), .B0(valid_mem[14]), .Y(n1237) );
  NAND2X1 U1052 ( .A(n1236), .B(n1235), .Y(n1083) );
  OAI21XL U1053 ( .A0(n1479), .A1(n855), .B0(valid_mem[13]), .Y(n1235) );
  NAND2X1 U1054 ( .A(n1234), .B(n1233), .Y(n1082) );
  OAI21XL U1055 ( .A0(n1476), .A1(n855), .B0(valid_mem[12]), .Y(n1233) );
  NAND2X1 U1056 ( .A(n1232), .B(n1231), .Y(n1081) );
  OAI21XL U1057 ( .A0(n1473), .A1(n855), .B0(valid_mem[11]), .Y(n1231) );
  NAND2X1 U1058 ( .A(n1228), .B(n1227), .Y(n1079) );
  OAI21XL U1059 ( .A0(n1467), .A1(n855), .B0(valid_mem[9]), .Y(n1227) );
  NAND2X1 U1060 ( .A(n1226), .B(n1225), .Y(n1078) );
  OAI21XL U1061 ( .A0(n1464), .A1(n855), .B0(valid_mem[8]), .Y(n1225) );
  NAND2X1 U1062 ( .A(n1222), .B(n1221), .Y(n1076) );
  OAI21XL U1063 ( .A0(n1458), .A1(n855), .B0(valid_mem[6]), .Y(n1221) );
  NAND2X1 U1064 ( .A(n1220), .B(n1219), .Y(n1075) );
  OAI21XL U1065 ( .A0(n1455), .A1(n855), .B0(valid_mem[5]), .Y(n1219) );
  NAND2X1 U1066 ( .A(n1218), .B(n1217), .Y(n1074) );
  OAI21XL U1067 ( .A0(n1452), .A1(n855), .B0(valid_mem[4]), .Y(n1217) );
  NAND2X1 U1068 ( .A(n1214), .B(n1213), .Y(n1072) );
  OAI21XL U1069 ( .A0(n1446), .A1(n855), .B0(valid_mem[2]), .Y(n1213) );
  NAND2X1 U1070 ( .A(n1224), .B(n1223), .Y(n1077) );
  OAI21XL U1071 ( .A0(n1461), .A1(n855), .B0(valid_mem[7]), .Y(n1223) );
  NAND2X1 U1072 ( .A(n1216), .B(n1215), .Y(n1073) );
  OAI21XL U1073 ( .A0(n1449), .A1(n855), .B0(valid_mem[3]), .Y(n1215) );
  NAND2X1 U1074 ( .A(n1212), .B(n1211), .Y(n1071) );
  OAI21XL U1075 ( .A0(n1443), .A1(n855), .B0(valid_mem[1]), .Y(n1211) );
  NAND2X1 U1076 ( .A(n1210), .B(n1209), .Y(n1070) );
  OAI21XL U1077 ( .A0(n1440), .A1(n855), .B0(valid_mem[0]), .Y(n1209) );
  NAND2X1 U1078 ( .A(n1389), .B(n1388), .Y(n1157) );
  OAI21XL U1079 ( .A0(n1461), .A1(n865), .B0(valid_mem[87]), .Y(n1388) );
endmodule


module LBP ( clk, reset, gray_addr, gray_req, gray_ready, gray_data, lbp_addr, 
        lbp_valid, lbp_data, finish );
  output [13:0] gray_addr;
  input [7:0] gray_data;
  output [13:0] lbp_addr;
  output [7:0] lbp_data;
  input clk, reset, gray_ready;
  output gray_req, lbp_valid, finish;
  wire   n265, line_buffer_1_valid, line_buffer_2_valid, \mask_data_out_3[1] ,
         \mask_data_out_6[1] , \mask_data_out_9[1] , n52, n54, n57, n58, n59,
         n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264;
  wire   [3:0] state;
  wire   [2:0] nstate;
  wire   [7:0] line_buffer_1_out;
  wire   [7:0] line_buffer_2_out;
  wire   [7:0] mask_data_out_1;
  wire   [7:0] mask_data_out_2;
  wire   [7:0] mask_data_out_4;
  wire   [7:0] mask_data_out_5;
  wire   [7:0] mask_data_out_7;
  wire   [7:0] mask_data_out_8;

  up_counter_WIDTH14_1 mem_addr_counter ( .clk(clk), .rst(n64), .clr(1'b0), 
        .count(gray_addr), .en_BAR(n79) );
  up_counter_WIDTH14_0 write_addr_counter ( .clk(clk), .rst(n64), .en(
        lbp_valid), .clr(1'b0), .count(lbp_addr) );
  line_buffer_1 line_buffer_1 ( .clk(clk), .rst(n64), .en(gray_req), .data_in(
        {n73, n72, n71, n70, n69, n68, n67, n66}), .data_out(line_buffer_1_out), .valid(line_buffer_1_valid) );
  line_buffer_0 line_buffer_2 ( .clk(clk), .rst(n64), .en(line_buffer_1_valid), 
        .data_in(line_buffer_1_out), .data_out(line_buffer_2_out), .valid(
        line_buffer_2_valid) );
  DFFRX1 lbp_valid_reg ( .D(n54), .CK(clk), .RN(n264), .Q(lbp_valid), .QN(n52)
         );
  EDFFX1 \mask_data_out_9_reg[1]  ( .D(mask_data_out_8[1]), .E(
        line_buffer_2_valid), .CK(clk), .Q(\mask_data_out_9[1] ) );
  EDFFX1 \mask_data_out_3_reg[1]  ( .D(mask_data_out_2[1]), .E(gray_req), .CK(
        clk), .Q(\mask_data_out_3[1] ) );
  EDFFX1 \mask_data_out_6_reg[1]  ( .D(mask_data_out_5[1]), .E(
        line_buffer_1_valid), .CK(clk), .Q(\mask_data_out_6[1] ) );
  EDFFX1 \mask_data_out_7_reg[1]  ( .D(line_buffer_2_out[1]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[1]) );
  EDFFX1 \mask_data_out_8_reg[1]  ( .D(mask_data_out_7[1]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[1]) );
  EDFFX1 \mask_data_out_1_reg[1]  ( .D(n67), .E(gray_req), .CK(clk), .Q(
        mask_data_out_1[1]) );
  EDFFX1 \mask_data_out_2_reg[1]  ( .D(mask_data_out_1[1]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[1]) );
  EDFFX1 \mask_data_out_4_reg[1]  ( .D(line_buffer_1_out[1]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[1]) );
  EDFFXL \mask_data_out_9_reg[7]  ( .D(mask_data_out_8[7]), .E(
        line_buffer_2_valid), .CK(clk), .QN(n252) );
  EDFFXL \mask_data_out_9_reg[6]  ( .D(mask_data_out_8[6]), .E(
        line_buffer_2_valid), .CK(clk), .QN(n261) );
  EDFFXL \mask_data_out_9_reg[5]  ( .D(mask_data_out_8[5]), .E(
        line_buffer_2_valid), .CK(clk), .Q(n196), .QN(n253) );
  EDFFXL \mask_data_out_9_reg[4]  ( .D(mask_data_out_8[4]), .E(
        line_buffer_2_valid), .CK(clk), .Q(n195) );
  EDFFXL \mask_data_out_9_reg[3]  ( .D(mask_data_out_8[3]), .E(
        line_buffer_2_valid), .CK(clk), .QN(n254) );
  EDFFXL \mask_data_out_9_reg[2]  ( .D(mask_data_out_8[2]), .E(
        line_buffer_2_valid), .CK(clk), .QN(n259) );
  EDFFXL \mask_data_out_9_reg[0]  ( .D(mask_data_out_8[0]), .E(
        line_buffer_2_valid), .CK(clk), .Q(n202), .QN(n258) );
  EDFFXL \mask_data_out_6_reg[7]  ( .D(mask_data_out_5[7]), .E(
        line_buffer_1_valid), .CK(clk), .Q(n57), .QN(n234) );
  EDFFXL \mask_data_out_6_reg[6]  ( .D(mask_data_out_5[6]), .E(
        line_buffer_1_valid), .CK(clk), .QN(n239) );
  EDFFXL \mask_data_out_6_reg[5]  ( .D(mask_data_out_5[5]), .E(
        line_buffer_1_valid), .CK(clk), .Q(n154), .QN(n235) );
  EDFFXL \mask_data_out_6_reg[4]  ( .D(mask_data_out_5[4]), .E(
        line_buffer_1_valid), .CK(clk), .Q(n153) );
  EDFFXL \mask_data_out_6_reg[3]  ( .D(mask_data_out_5[3]), .E(
        line_buffer_1_valid), .CK(clk), .QN(n236) );
  EDFFXL \mask_data_out_6_reg[2]  ( .D(mask_data_out_5[2]), .E(
        line_buffer_1_valid), .CK(clk), .QN(n238) );
  EDFFXL \mask_data_out_6_reg[0]  ( .D(mask_data_out_5[0]), .E(
        line_buffer_1_valid), .CK(clk), .Q(n160), .QN(n237) );
  EDFFXL \mask_data_out_3_reg[7]  ( .D(mask_data_out_2[7]), .E(gray_req), .CK(
        clk), .Q(n59), .QN(n222) );
  EDFFXL \mask_data_out_3_reg[6]  ( .D(mask_data_out_2[6]), .E(gray_req), .CK(
        clk), .QN(n227) );
  EDFFXL \mask_data_out_3_reg[5]  ( .D(mask_data_out_2[5]), .E(gray_req), .CK(
        clk), .Q(n125), .QN(n223) );
  EDFFXL \mask_data_out_3_reg[4]  ( .D(mask_data_out_2[4]), .E(gray_req), .CK(
        clk), .Q(n124) );
  EDFFXL \mask_data_out_3_reg[3]  ( .D(mask_data_out_2[3]), .E(gray_req), .CK(
        clk), .QN(n224) );
  EDFFXL \mask_data_out_3_reg[2]  ( .D(mask_data_out_2[2]), .E(gray_req), .CK(
        clk), .QN(n226) );
  EDFFXL \mask_data_out_3_reg[0]  ( .D(mask_data_out_2[0]), .E(gray_req), .CK(
        clk), .Q(n131), .QN(n225) );
  EDFFXL \mask_data_out_8_reg[7]  ( .D(mask_data_out_7[7]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[7]), .QN(n246) );
  EDFFXL \mask_data_out_8_reg[6]  ( .D(mask_data_out_7[6]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[6]), .QN(n251) );
  EDFFXL \mask_data_out_8_reg[5]  ( .D(mask_data_out_7[5]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[5]), .QN(n247) );
  EDFFXL \mask_data_out_8_reg[4]  ( .D(mask_data_out_7[4]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[4]) );
  EDFFXL \mask_data_out_8_reg[3]  ( .D(mask_data_out_7[3]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[3]), .QN(n248) );
  EDFFXL \mask_data_out_8_reg[2]  ( .D(mask_data_out_7[2]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[2]), .QN(n250) );
  EDFFXL \mask_data_out_8_reg[0]  ( .D(mask_data_out_7[0]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_8[0]), .QN(n249) );
  EDFFXL \mask_data_out_7_reg[7]  ( .D(line_buffer_2_out[7]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[7]), .QN(n240) );
  EDFFXL \mask_data_out_7_reg[6]  ( .D(line_buffer_2_out[6]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[6]), .QN(n245) );
  EDFFXL \mask_data_out_7_reg[5]  ( .D(line_buffer_2_out[5]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[5]), .QN(n241) );
  EDFFXL \mask_data_out_7_reg[4]  ( .D(line_buffer_2_out[4]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[4]) );
  EDFFXL \mask_data_out_7_reg[3]  ( .D(line_buffer_2_out[3]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[3]), .QN(n242) );
  EDFFXL \mask_data_out_7_reg[2]  ( .D(line_buffer_2_out[2]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[2]), .QN(n244) );
  EDFFXL \mask_data_out_7_reg[0]  ( .D(line_buffer_2_out[0]), .E(
        line_buffer_2_valid), .CK(clk), .Q(mask_data_out_7[0]), .QN(n243) );
  EDFFXL \mask_data_out_5_reg[0]  ( .D(mask_data_out_4[0]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[0]), .QN(n255) );
  EDFFXL \mask_data_out_4_reg[7]  ( .D(line_buffer_1_out[7]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[7]), .QN(n228) );
  EDFFXL \mask_data_out_4_reg[6]  ( .D(line_buffer_1_out[6]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[6]), .QN(n233) );
  EDFFXL \mask_data_out_4_reg[5]  ( .D(line_buffer_1_out[5]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[5]), .QN(n229) );
  EDFFXL \mask_data_out_4_reg[4]  ( .D(line_buffer_1_out[4]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[4]) );
  EDFFXL \mask_data_out_4_reg[3]  ( .D(line_buffer_1_out[3]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[3]), .QN(n230) );
  EDFFXL \mask_data_out_4_reg[2]  ( .D(line_buffer_1_out[2]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[2]), .QN(n232) );
  EDFFXL \mask_data_out_4_reg[0]  ( .D(line_buffer_1_out[0]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_4[0]), .QN(n231) );
  EDFFXL \mask_data_out_2_reg[7]  ( .D(mask_data_out_1[7]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[7]), .QN(n216) );
  EDFFXL \mask_data_out_2_reg[6]  ( .D(mask_data_out_1[6]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[6]), .QN(n221) );
  EDFFXL \mask_data_out_2_reg[5]  ( .D(mask_data_out_1[5]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[5]), .QN(n217) );
  EDFFXL \mask_data_out_2_reg[4]  ( .D(mask_data_out_1[4]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[4]) );
  EDFFXL \mask_data_out_2_reg[3]  ( .D(mask_data_out_1[3]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[3]), .QN(n218) );
  EDFFXL \mask_data_out_2_reg[2]  ( .D(mask_data_out_1[2]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[2]), .QN(n220) );
  EDFFXL \mask_data_out_2_reg[0]  ( .D(mask_data_out_1[0]), .E(gray_req), .CK(
        clk), .Q(mask_data_out_2[0]), .QN(n219) );
  EDFFXL \mask_data_out_1_reg[7]  ( .D(gray_data[7]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[7]), .QN(n210) );
  EDFFXL \mask_data_out_1_reg[6]  ( .D(gray_data[6]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[6]), .QN(n215) );
  EDFFXL \mask_data_out_1_reg[5]  ( .D(gray_data[5]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[5]), .QN(n211) );
  EDFFXL \mask_data_out_1_reg[4]  ( .D(gray_data[4]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[4]), .QN(n61) );
  EDFFXL \mask_data_out_1_reg[3]  ( .D(gray_data[3]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[3]), .QN(n212) );
  EDFFXL \mask_data_out_1_reg[2]  ( .D(gray_data[2]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[2]), .QN(n214) );
  EDFFXL \mask_data_out_1_reg[0]  ( .D(gray_data[0]), .E(gray_req), .CK(clk), 
        .Q(mask_data_out_1[0]), .QN(n213) );
  DFFRX1 \state_reg[2]  ( .D(nstate[2]), .CK(clk), .RN(n264), .Q(state[2]), 
        .QN(n60) );
  DFFRX1 \state_reg[1]  ( .D(nstate[1]), .CK(clk), .RN(n264), .Q(state[1]), 
        .QN(n58) );
  DFFRX1 \state_reg[0]  ( .D(nstate[0]), .CK(clk), .RN(n264), .Q(state[0]), 
        .QN(n82) );
  EDFFX4 \mask_data_out_5_reg[6]  ( .D(mask_data_out_4[6]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[6]) );
  EDFFX4 \mask_data_out_5_reg[3]  ( .D(mask_data_out_4[3]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[3]) );
  EDFFX4 \mask_data_out_5_reg[2]  ( .D(mask_data_out_4[2]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[2]), .QN(n260) );
  EDFFX2 \mask_data_out_5_reg[1]  ( .D(mask_data_out_4[1]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[1]), .QN(n257) );
  EDFFX2 \mask_data_out_5_reg[7]  ( .D(mask_data_out_4[7]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[7]), .QN(n256) );
  EDFFX2 \mask_data_out_5_reg[5]  ( .D(mask_data_out_4[5]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[5]), .QN(n262) );
  EDFFX2 \mask_data_out_5_reg[4]  ( .D(mask_data_out_4[4]), .E(
        line_buffer_1_valid), .CK(clk), .Q(mask_data_out_5[4]), .QN(n263) );
  NOR2X1 U52 ( .A(n57), .B(n256), .Y(n146) );
  NOR2X1 U53 ( .A(mask_data_out_4[7]), .B(n256), .Y(n133) );
  NAND3X1 U54 ( .A(n58), .B(n82), .C(state[2]), .Y(n81) );
  NOR2X1 U55 ( .A(n59), .B(n256), .Y(n117) );
  NOR2X1 U56 ( .A(mask_data_out_2[7]), .B(n256), .Y(n104) );
  NAND4X1 U57 ( .A(n60), .B(state[1]), .C(gray_ready), .D(n82), .Y(n80) );
  NAND2X1 U58 ( .A(mask_data_out_5[0]), .B(mask_data_out_5[1]), .Y(n102) );
  AOI22X1 U59 ( .A0(mask_data_out_5[6]), .A1(n215), .B0(mask_data_out_5[4]), 
        .B1(n61), .Y(n92) );
  NAND3X1 U60 ( .A(n77), .B(n76), .C(n52), .Y(n54) );
  INVXL U61 ( .A(n265), .Y(n62) );
  INVX4 U62 ( .A(n62), .Y(gray_req) );
  AND2XL U63 ( .A(n200), .B(n260), .Y(n199) );
  AOI2BB1XL U64 ( .A0N(n200), .A1N(n260), .B0(n259), .Y(n198) );
  AND2XL U65 ( .A(n185), .B(n260), .Y(n184) );
  AOI2BB1XL U66 ( .A0N(n185), .A1N(n260), .B0(n250), .Y(n183) );
  AND2XL U67 ( .A(n172), .B(n260), .Y(n171) );
  AOI2BB1XL U68 ( .A0N(n172), .A1N(n260), .B0(n244), .Y(n170) );
  AND2XL U69 ( .A(n158), .B(n260), .Y(n157) );
  AOI2BB1XL U70 ( .A0N(n158), .A1N(n260), .B0(n238), .Y(n156) );
  AND2XL U71 ( .A(n143), .B(n260), .Y(n142) );
  AOI2BB1XL U72 ( .A0N(n143), .A1N(n260), .B0(n232), .Y(n141) );
  AND2XL U73 ( .A(n129), .B(n260), .Y(n128) );
  AOI2BB1XL U74 ( .A0N(n129), .A1N(n260), .B0(n226), .Y(n127) );
  AND2XL U75 ( .A(n114), .B(n260), .Y(n113) );
  AOI2BB1XL U76 ( .A0N(n114), .A1N(n260), .B0(n220), .Y(n112) );
  AND2XL U77 ( .A(n99), .B(n260), .Y(n98) );
  AOI2BB1XL U78 ( .A0N(n99), .A1N(n260), .B0(n214), .Y(n97) );
  OAI211XL U79 ( .A0(n258), .A1(mask_data_out_5[1]), .B0(n201), .C0(n101), .Y(
        n200) );
  OAI211XL U80 ( .A0(n249), .A1(mask_data_out_5[1]), .B0(n186), .C0(n101), .Y(
        n185) );
  OAI211XL U81 ( .A0(n243), .A1(mask_data_out_5[1]), .B0(n173), .C0(n101), .Y(
        n172) );
  OAI211XL U82 ( .A0(n237), .A1(mask_data_out_5[1]), .B0(n159), .C0(n101), .Y(
        n158) );
  OAI211XL U83 ( .A0(n231), .A1(mask_data_out_5[1]), .B0(n144), .C0(n101), .Y(
        n143) );
  OAI211XL U84 ( .A0(n225), .A1(mask_data_out_5[1]), .B0(n130), .C0(n101), .Y(
        n129) );
  OAI211XL U85 ( .A0(n219), .A1(mask_data_out_5[1]), .B0(n115), .C0(n101), .Y(
        n114) );
  OAI211XL U86 ( .A0(n213), .A1(mask_data_out_5[1]), .B0(n100), .C0(n101), .Y(
        n99) );
  OAI32XL U87 ( .A0(n65), .A1(n187), .A2(n188), .B0(n252), .B1(n89), .Y(
        lbp_data[0]) );
  AOI2BB2XL U88 ( .B0(mask_data_out_5[6]), .B1(n261), .A0N(n263), .A1N(n195), 
        .Y(n191) );
  OAI32XL U89 ( .A0(n65), .A1(n174), .A2(n175), .B0(n246), .B1(n89), .Y(
        lbp_data[1]) );
  AOI2BB2XL U90 ( .B0(mask_data_out_5[6]), .B1(n251), .A0N(n263), .A1N(
        mask_data_out_8[4]), .Y(n178) );
  OAI32XL U91 ( .A0(n65), .A1(n161), .A2(n162), .B0(n240), .B1(n89), .Y(
        lbp_data[2]) );
  AOI2BB2XL U92 ( .B0(mask_data_out_5[6]), .B1(n245), .A0N(n263), .A1N(
        mask_data_out_7[4]), .Y(n165) );
  OAI32XL U93 ( .A0(n65), .A1(n145), .A2(n146), .B0(n234), .B1(n89), .Y(
        lbp_data[3]) );
  AOI2BB2XL U94 ( .B0(mask_data_out_5[6]), .B1(n239), .A0N(n263), .A1N(n153), 
        .Y(n149) );
  OAI32XL U95 ( .A0(n65), .A1(n132), .A2(n133), .B0(n228), .B1(n89), .Y(
        lbp_data[4]) );
  AOI2BB2XL U96 ( .B0(mask_data_out_5[6]), .B1(n233), .A0N(n263), .A1N(
        mask_data_out_4[4]), .Y(n136) );
  OAI32XL U97 ( .A0(n65), .A1(n116), .A2(n117), .B0(n222), .B1(n89), .Y(
        lbp_data[5]) );
  AOI2BB2XL U98 ( .B0(mask_data_out_5[6]), .B1(n227), .A0N(n263), .A1N(n124), 
        .Y(n120) );
  OAI32XL U99 ( .A0(n65), .A1(n103), .A2(n104), .B0(n216), .B1(n89), .Y(
        lbp_data[6]) );
  AOI2BB2XL U100 ( .B0(mask_data_out_5[6]), .B1(n221), .A0N(n263), .A1N(
        mask_data_out_2[4]), .Y(n107) );
  OAI32XL U101 ( .A0(n65), .A1(n87), .A2(n88), .B0(n210), .B1(n89), .Y(
        lbp_data[7]) );
  AOI32XL U102 ( .A0(n263), .A1(mask_data_out_8[4]), .A2(n176), .B0(
        mask_data_out_8[5]), .B1(n262), .Y(n181) );
  AOI32XL U103 ( .A0(n263), .A1(mask_data_out_7[4]), .A2(n163), .B0(
        mask_data_out_7[5]), .B1(n262), .Y(n168) );
  AOI32XL U104 ( .A0(n263), .A1(n153), .A2(n147), .B0(n154), .B1(n262), .Y(
        n152) );
  AOI32XL U105 ( .A0(n263), .A1(mask_data_out_4[4]), .A2(n134), .B0(
        mask_data_out_4[5]), .B1(n262), .Y(n139) );
  AOI32XL U106 ( .A0(n263), .A1(n124), .A2(n118), .B0(n125), .B1(n262), .Y(
        n123) );
  AOI32XL U107 ( .A0(n263), .A1(mask_data_out_2[4]), .A2(n105), .B0(
        mask_data_out_2[5]), .B1(n262), .Y(n110) );
  AOI32XL U108 ( .A0(n263), .A1(mask_data_out_1[4]), .A2(n90), .B0(
        mask_data_out_1[5]), .B1(n262), .Y(n95) );
  AOI32XL U109 ( .A0(n263), .A1(n195), .A2(n189), .B0(n196), .B1(n262), .Y(
        n194) );
  NAND2XL U110 ( .A(n253), .B(mask_data_out_5[5]), .Y(n189) );
  NAND2XL U111 ( .A(n247), .B(mask_data_out_5[5]), .Y(n176) );
  NAND2XL U112 ( .A(n241), .B(mask_data_out_5[5]), .Y(n163) );
  NAND2XL U113 ( .A(n235), .B(mask_data_out_5[5]), .Y(n147) );
  NAND2XL U114 ( .A(n229), .B(mask_data_out_5[5]), .Y(n134) );
  NAND2XL U115 ( .A(n223), .B(mask_data_out_5[5]), .Y(n118) );
  NAND2XL U116 ( .A(n217), .B(mask_data_out_5[5]), .Y(n105) );
  NAND2XL U117 ( .A(n211), .B(mask_data_out_5[5]), .Y(n90) );
  CLKBUFX3 U118 ( .A(n86), .Y(n65) );
  OAI221XL U119 ( .A0(n203), .A1(n204), .B0(n205), .B1(n206), .C0(n207), .Y(
        n86) );
  CLKBUFX3 U120 ( .A(gray_data[0]), .Y(n66) );
  CLKBUFX3 U121 ( .A(gray_data[1]), .Y(n67) );
  CLKBUFX3 U122 ( .A(gray_data[2]), .Y(n68) );
  CLKBUFX3 U123 ( .A(gray_data[3]), .Y(n69) );
  CLKBUFX3 U124 ( .A(gray_data[4]), .Y(n70) );
  CLKBUFX3 U125 ( .A(gray_data[5]), .Y(n71) );
  CLKBUFX3 U126 ( .A(gray_data[6]), .Y(n72) );
  CLKBUFX3 U127 ( .A(gray_data[7]), .Y(n73) );
  CLKBUFX3 U128 ( .A(reset), .Y(n64) );
  OR4X1 U129 ( .A(gray_addr[4]), .B(gray_addr[3]), .C(gray_addr[6]), .D(
        gray_addr[5]), .Y(n74) );
  OR4X1 U130 ( .A(gray_addr[2]), .B(gray_addr[1]), .C(gray_addr[0]), .D(n74), 
        .Y(n75) );
  AOI211X1 U131 ( .A0(gray_addr[7]), .A1(n75), .B0(gray_addr[11]), .C0(
        gray_addr[10]), .Y(n77) );
  NOR4X1 U132 ( .A(gray_addr[9]), .B(gray_addr[8]), .C(gray_addr[13]), .D(
        gray_addr[12]), .Y(n76) );
  OAI211X1 U133 ( .A0(n78), .A1(n79), .B0(n80), .C0(n81), .Y(nstate[2]) );
  OAI2BB2XL U134 ( .B0(n78), .B1(n79), .A0N(n83), .A1N(n82), .Y(nstate[1]) );
  OAI21XL U135 ( .A0(state[2]), .A1(gray_ready), .B0(state[1]), .Y(n83) );
  AND2X1 U136 ( .A(n84), .B(n85), .Y(n78) );
  OR2X1 U137 ( .A(finish), .B(n265), .Y(nstate[0]) );
  CLKINVX1 U138 ( .A(n64), .Y(n264) );
  NOR2BX1 U139 ( .AN(n210), .B(n256), .Y(n88) );
  AOI32X1 U140 ( .A0(n90), .A1(n91), .A2(n92), .B0(n93), .B1(n94), .Y(n87) );
  OAI21XL U141 ( .A0(n95), .A1(mask_data_out_5[6]), .B0(n215), .Y(n94) );
  NAND2X1 U142 ( .A(n95), .B(mask_data_out_5[6]), .Y(n93) );
  OAI21XL U143 ( .A0(n212), .A1(mask_data_out_5[3]), .B0(n96), .Y(n91) );
  OAI2BB2XL U144 ( .B0(n97), .B1(n98), .A0N(mask_data_out_5[3]), .A1N(n212), 
        .Y(n96) );
  OAI21XL U145 ( .A0(n102), .A1(mask_data_out_1[0]), .B0(mask_data_out_1[1]), 
        .Y(n100) );
  AOI32X1 U146 ( .A0(n105), .A1(n106), .A2(n107), .B0(n108), .B1(n109), .Y(
        n103) );
  OAI21XL U147 ( .A0(n110), .A1(mask_data_out_5[6]), .B0(n221), .Y(n109) );
  NAND2X1 U148 ( .A(n110), .B(mask_data_out_5[6]), .Y(n108) );
  OAI21XL U149 ( .A0(n218), .A1(mask_data_out_5[3]), .B0(n111), .Y(n106) );
  OAI2BB2XL U150 ( .B0(n112), .B1(n113), .A0N(mask_data_out_5[3]), .A1N(n218), 
        .Y(n111) );
  OAI21XL U151 ( .A0(n102), .A1(mask_data_out_2[0]), .B0(mask_data_out_2[1]), 
        .Y(n115) );
  AOI32X1 U152 ( .A0(n118), .A1(n119), .A2(n120), .B0(n121), .B1(n122), .Y(
        n116) );
  OAI21XL U153 ( .A0(n123), .A1(mask_data_out_5[6]), .B0(n227), .Y(n122) );
  NAND2X1 U154 ( .A(n123), .B(mask_data_out_5[6]), .Y(n121) );
  OAI21XL U155 ( .A0(n224), .A1(mask_data_out_5[3]), .B0(n126), .Y(n119) );
  OAI2BB2XL U156 ( .B0(n127), .B1(n128), .A0N(mask_data_out_5[3]), .A1N(n224), 
        .Y(n126) );
  OAI21XL U157 ( .A0(n102), .A1(n131), .B0(\mask_data_out_3[1] ), .Y(n130) );
  AOI32X1 U158 ( .A0(n134), .A1(n135), .A2(n136), .B0(n137), .B1(n138), .Y(
        n132) );
  OAI21XL U159 ( .A0(n139), .A1(mask_data_out_5[6]), .B0(n233), .Y(n138) );
  NAND2X1 U160 ( .A(n139), .B(mask_data_out_5[6]), .Y(n137) );
  OAI21XL U161 ( .A0(n230), .A1(mask_data_out_5[3]), .B0(n140), .Y(n135) );
  OAI2BB2XL U162 ( .B0(n141), .B1(n142), .A0N(mask_data_out_5[3]), .A1N(n230), 
        .Y(n140) );
  OAI21XL U163 ( .A0(n102), .A1(mask_data_out_4[0]), .B0(mask_data_out_4[1]), 
        .Y(n144) );
  AOI32X1 U164 ( .A0(n147), .A1(n148), .A2(n149), .B0(n150), .B1(n151), .Y(
        n145) );
  OAI21XL U165 ( .A0(n152), .A1(mask_data_out_5[6]), .B0(n239), .Y(n151) );
  NAND2X1 U166 ( .A(n152), .B(mask_data_out_5[6]), .Y(n150) );
  OAI21XL U167 ( .A0(n236), .A1(mask_data_out_5[3]), .B0(n155), .Y(n148) );
  OAI2BB2XL U168 ( .B0(n156), .B1(n157), .A0N(mask_data_out_5[3]), .A1N(n236), 
        .Y(n155) );
  OAI21XL U169 ( .A0(n102), .A1(n160), .B0(\mask_data_out_6[1] ), .Y(n159) );
  NOR2BX1 U170 ( .AN(n240), .B(n256), .Y(n162) );
  AOI32X1 U171 ( .A0(n163), .A1(n164), .A2(n165), .B0(n166), .B1(n167), .Y(
        n161) );
  OAI21XL U172 ( .A0(n168), .A1(mask_data_out_5[6]), .B0(n245), .Y(n167) );
  NAND2X1 U173 ( .A(n168), .B(mask_data_out_5[6]), .Y(n166) );
  OAI21XL U174 ( .A0(n242), .A1(mask_data_out_5[3]), .B0(n169), .Y(n164) );
  OAI2BB2XL U175 ( .B0(n170), .B1(n171), .A0N(mask_data_out_5[3]), .A1N(n242), 
        .Y(n169) );
  OAI21XL U176 ( .A0(n102), .A1(mask_data_out_7[0]), .B0(mask_data_out_7[1]), 
        .Y(n173) );
  NOR2BX1 U177 ( .AN(n246), .B(n256), .Y(n175) );
  AOI32X1 U178 ( .A0(n176), .A1(n177), .A2(n178), .B0(n179), .B1(n180), .Y(
        n174) );
  OAI21XL U179 ( .A0(n181), .A1(mask_data_out_5[6]), .B0(n251), .Y(n180) );
  NAND2X1 U180 ( .A(n181), .B(mask_data_out_5[6]), .Y(n179) );
  OAI21XL U181 ( .A0(n248), .A1(mask_data_out_5[3]), .B0(n182), .Y(n177) );
  OAI2BB2XL U182 ( .B0(n183), .B1(n184), .A0N(mask_data_out_5[3]), .A1N(n248), 
        .Y(n182) );
  OAI21XL U183 ( .A0(n102), .A1(mask_data_out_8[0]), .B0(mask_data_out_8[1]), 
        .Y(n186) );
  NAND2BX1 U184 ( .AN(n65), .B(n256), .Y(n89) );
  NOR2BX1 U185 ( .AN(n252), .B(n256), .Y(n188) );
  AOI32X1 U186 ( .A0(n189), .A1(n190), .A2(n191), .B0(n192), .B1(n193), .Y(
        n187) );
  OAI21XL U187 ( .A0(n194), .A1(n261), .B0(mask_data_out_5[6]), .Y(n193) );
  NAND2X1 U188 ( .A(n194), .B(n261), .Y(n192) );
  OAI21XL U189 ( .A0(n254), .A1(mask_data_out_5[3]), .B0(n197), .Y(n190) );
  OAI2BB2XL U190 ( .B0(n198), .B1(n199), .A0N(mask_data_out_5[3]), .A1N(n254), 
        .Y(n197) );
  NAND2X1 U191 ( .A(n255), .B(n257), .Y(n101) );
  OAI21XL U192 ( .A0(n102), .A1(n202), .B0(\mask_data_out_9[1] ), .Y(n201) );
  NOR2X1 U193 ( .A(n84), .B(n85), .Y(n207) );
  AND4X1 U194 ( .A(lbp_addr[5]), .B(lbp_addr[4]), .C(lbp_addr[6]), .D(n208), 
        .Y(n85) );
  AND4X1 U195 ( .A(lbp_addr[0]), .B(lbp_addr[1]), .C(lbp_addr[2]), .D(
        lbp_addr[3]), .Y(n208) );
  AND4X1 U196 ( .A(lbp_addr[8]), .B(lbp_addr[7]), .C(lbp_addr[9]), .D(n209), 
        .Y(n84) );
  AND4X1 U197 ( .A(lbp_addr[10]), .B(lbp_addr[11]), .C(lbp_addr[12]), .D(
        lbp_addr[13]), .Y(n209) );
  OR3X1 U198 ( .A(lbp_addr[11]), .B(lbp_addr[12]), .C(lbp_addr[10]), .Y(n206)
         );
  OR4X1 U199 ( .A(lbp_addr[13]), .B(lbp_addr[7]), .C(lbp_addr[8]), .D(
        lbp_addr[9]), .Y(n205) );
  OR3X1 U200 ( .A(lbp_addr[1]), .B(lbp_addr[2]), .C(lbp_addr[0]), .Y(n204) );
  OR4X1 U201 ( .A(lbp_addr[3]), .B(lbp_addr[4]), .C(lbp_addr[5]), .D(
        lbp_addr[6]), .Y(n203) );
  NAND2X1 U202 ( .A(n79), .B(n81), .Y(n265) );
  NAND3X1 U203 ( .A(state[1]), .B(state[2]), .C(state[0]), .Y(n79) );
  NOR3X1 U204 ( .A(state[1]), .B(state[2]), .C(n82), .Y(finish) );
endmodule

